`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company:
// Engineer:
//
// Create Date: 24.01.2020 18:13:04
// Design Name:
// Module Name: test
// Project Name:
// Target Devices:
// Tool Versions:
// Description:
//
// Dependencies:
//
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
//
//////////////////////////////////////////////////////////////////////////////////


module simulation();
reg clk,reset;
//reg [5:0]in;
reg [31:0]value1,value2;
wire [63:0]op1,op2;
//wire vaouten;
integer handle1;
//topmod m1 (clk,reset,value1,value2,op1,op2);
wire [9:0] addrext;
 wire valid;
 wire zeros;
 wire done;
topmod m1(clk,reset,value1,value2,addrext,valid,zeros,op1,op2,done);
/* 
input clk;
input reset;
input[31:0] input1;
input [31:0]input2;
output wire [63:0] op1;
output wire [63:0] op2;
output 
 */


initial begin
reset=0;
value1=0;
value2=0;
clk=0;
end

initial
begin
#70 clk=0;
forever #200 clk=~clk;
end
initial begin
#50 reset=0;
end
initial begin
#450 reset=0;
#400 reset=1;
end
/*
//alpha_post rgr (clk,reset,temp,vaout,vaouten);
initial
begin

 handle1 = $fopen("file1.out");

end

always@(posedge clk) begin
if(vaouten==0) begin
end
else if(vaouten==1) begin 
$fdisplay(handle1,"%d",vaout);
end
end
*/
//initial begin
//#10000000 $finish;
//end
/*
initial
clk=1'b0;
initial
reset=0;

initial
#110 reset=1;
initial
#120 reset=0;
*/
initial
begin 
//value
#450 value1=32'd1;value2=32'd1;
#1747200 value1=32'd1;value2=32'd1;
//column
#400 value1=32'd1;value2=32'd4;
#400 value1=32'd5;value2=32'd6;
#400 value1=32'd8;value2=32'd14;
#400 value1=32'd15;value2=32'd16;
#400 value1=32'd20;value2=32'd22;
#400 value1=32'd106;value2=32'd107;
#400 value1=32'd110;value2=32'd112;
#400 value1=32'd0;value2=32'd4;
#400 value1=32'd5;value2=32'd7;
#400 value1=32'd9;value2=32'd27;
#400 value1=32'd28;value2=32'd32;
#400 value1=32'd34;value2=32'd105;
#400 value1=32'd118;value2=32'd119;
#400 value1=32'd122;value2=32'd124;
#400 value1=32'd3;value2=32'd4;
#400 value1=32'd10;value2=32'd12;
#400 value1=32'd27;value2=32'd39;
#400 value1=32'd43;value2=32'd45;
#400 value1=32'd106;value2=32'd130;
#400 value1=32'd133;value2=32'd135;
#400 value1=32'd2;value2=32'd5;
#400 value1=32'd11;value2=32'd13;
#400 value1=32'd28;value2=32'd39;
#400 value1=32'd53;value2=32'd55;
#400 value1=32'd107;value2=32'd130;
#400 value1=32'd143;value2=32'd145;
#400 value1=32'd0;value2=32'd1;
#400 value1=32'd2;value2=32'd5;
#400 value1=32'd10;value2=32'd12;
#400 value1=32'd29;value2=32'd40;
#400 value1=32'd50;value2=32'd62;
#400 value1=32'd64;value2=32'd108;
#400 value1=32'd131;value2=32'd141;
#400 value1=32'd152;value2=32'd154;
#400 value1=32'd0;value2=32'd1;
#400 value1=32'd3;value2=32'd4;
#400 value1=32'd11;value2=32'd13;
#400 value1=32'd30;value2=32'd41;
#400 value1=32'd51;value2=32'd70;
#400 value1=32'd72;value2=32'd109;
#400 value1=32'd132;value2=32'd142;
#400 value1=32'd160;value2=32'd162;
#400 value1=32'd0;value2=32'd7;
#400 value1=32'd8;value2=32'd10;
#400 value1=32'd11;value2=32'd31;
#400 value1=32'd42;value2=32'd52;
#400 value1=32'd77;value2=32'd79;
#400 value1=32'd110;value2=32'd133;
#400 value1=32'd143;value2=32'd169;
#400 value1=32'd1;value2=32'd6;
#400 value1=32'd9;value2=32'd10;
#400 value1=32'd11;value2=32'd32;
#400 value1=32'd43;value2=32'd53;
#400 value1=32'd85;value2=32'd111;
#400 value1=32'd134;value2=32'd144;
#400 value1=32'd168;value2=32'd175;
#400 value1=32'd0;value2=32'd6;
#400 value1=32'd9;value2=32'd12;
#400 value1=32'd13;value2=32'd33;
#400 value1=32'd44;value2=32'd54;
#400 value1=32'd84;value2=32'd90;
#400 value1=32'd112;value2=32'd135;
#400 value1=32'd145;value2=32'd169;
#400 value1=32'd1;value2=32'd7;
#400 value1=32'd8;value2=32'd12;
#400 value1=32'd13;value2=32'd34;
#400 value1=32'd45;value2=32'd55;
#400 value1=32'd85;value2=32'd113;
#400 value1=32'd136;value2=32'd146;
#400 value1=32'd170;value2=32'd181;
#400 value1=32'd2;value2=32'd4;
#400 value1=32'd6;value2=32'd7;
#400 value1=32'd11;value2=32'd12;
#400 value1=32'd35;value2=32'd46;
#400 value1=32'd56;value2=32'd86;
#400 value1=32'd95;value2=32'd114;
#400 value1=32'd137;value2=32'd147;
#400 value1=32'd171;value2=32'd182;
#400 value1=32'd3;value2=32'd5;
#400 value1=32'd6;value2=32'd7;
#400 value1=32'd10;value2=32'd13;
#400 value1=32'd36;value2=32'd47;
#400 value1=32'd57;value2=32'd87;
#400 value1=32'd96;value2=32'd115;
#400 value1=32'd138;value2=32'd148;
#400 value1=32'd172;value2=32'd183;
#400 value1=32'd2;value2=32'd4;
#400 value1=32'd8;value2=32'd9;
#400 value1=32'd10;value2=32'd13;
#400 value1=32'd37;value2=32'd48;
#400 value1=32'd58;value2=32'd88;
#400 value1=32'd97;value2=32'd116;
#400 value1=32'd139;value2=32'd149;
#400 value1=32'd173;value2=32'd184;
#400 value1=32'd3;value2=32'd5;
#400 value1=32'd8;value2=32'd9;
#400 value1=32'd11;value2=32'd12;
#400 value1=32'd38;value2=32'd49;
#400 value1=32'd59;value2=32'd89;
#400 value1=32'd98;value2=32'd117;
#400 value1=32'd140;value2=32'd150;
#400 value1=32'd174;value2=32'd185;
#400 value1=32'd0;value2=32'd17;
#400 value1=32'd18;value2=32'd20;
#400 value1=32'd22;value2=32'd29;
#400 value1=32'd30;value2=32'd31;
#400 value1=32'd33;value2=32'd105;
#400 value1=32'd196;value2=32'd197;
#400 value1=32'd200;value2=32'd202;
#400 value1=32'd0;value2=32'd16;
#400 value1=32'd17;value2=32'd23;
#400 value1=32'd25;value2=32'd27;
#400 value1=32'd40;value2=32'd41;
#400 value1=32'd42;value2=32'd44;
#400 value1=32'd106;value2=32'd208;
#400 value1=32'd211;value2=32'd213;
#400 value1=32'd0;value2=32'd15;
#400 value1=32'd18;value2=32'd24;
#400 value1=32'd26;value2=32'd28;
#400 value1=32'd50;value2=32'd51;
#400 value1=32'd52;value2=32'd54;
#400 value1=32'd107;value2=32'd208;
#400 value1=32'd221;value2=32'd223;
#400 value1=32'd14;value2=32'd15;
#400 value1=32'd18;value2=32'd23;
#400 value1=32'd25;value2=32'd29;
#400 value1=32'd60;value2=32'd61;
#400 value1=32'd63;value2=32'd108;
#400 value1=32'd209;value2=32'd219;
#400 value1=32'd230;value2=32'd232;
#400 value1=32'd14;value2=32'd16;
#400 value1=32'd17;value2=32'd24;
#400 value1=32'd26;value2=32'd30;
#400 value1=32'd60;value2=32'd69;
#400 value1=32'd71;value2=32'd109;
#400 value1=32'd210;value2=32'd220;
#400 value1=32'd238;value2=32'd240;
#400 value1=32'd20;value2=32'd21;
#400 value1=32'd23;value2=32'd24;
#400 value1=32'd31;value2=32'd61;
#400 value1=32'd69;value2=32'd78;
#400 value1=32'd110;value2=32'd211;
#400 value1=32'd221;value2=32'd247;
#400 value1=32'd0;value2=32'd14;
#400 value1=32'd19;value2=32'd22;
#400 value1=32'd23;value2=32'd24;
#400 value1=32'd32;value2=32'd62;
#400 value1=32'd70;value2=32'd77;
#400 value1=32'd84;value2=32'd111;
#400 value1=32'd212;value2=32'd222;
#400 value1=32'd246;value2=32'd253;
#400 value1=32'd19;value2=32'd22;
#400 value1=32'd25;value2=32'd26;
#400 value1=32'd33;value2=32'd63;
#400 value1=32'd71;value2=32'd78;
#400 value1=32'd112;value2=32'd213;
#400 value1=32'd223;value2=32'd247;
#400 value1=32'd0;value2=32'd14;
#400 value1=32'd20;value2=32'd21;
#400 value1=32'd25;value2=32'd26;
#400 value1=32'd34;value2=32'd64;
#400 value1=32'd72;value2=32'd79;
#400 value1=32'd90;value2=32'd113;
#400 value1=32'd214;value2=32'd224;
#400 value1=32'd248;value2=32'd259;
#400 value1=32'd15;value2=32'd17;
#400 value1=32'd19;value2=32'd20;
#400 value1=32'd24;value2=32'd25;
#400 value1=32'd35;value2=32'd65;
#400 value1=32'd73;value2=32'd80;
#400 value1=32'd91;value2=32'd114;
#400 value1=32'd215;value2=32'd225;
#400 value1=32'd249;value2=32'd260;
#400 value1=32'd16;value2=32'd18;
#400 value1=32'd19;value2=32'd20;
#400 value1=32'd23;value2=32'd26;
#400 value1=32'd36;value2=32'd66;
#400 value1=32'd74;value2=32'd81;
#400 value1=32'd92;value2=32'd115;
#400 value1=32'd216;value2=32'd226;
#400 value1=32'd250;value2=32'd261;
#400 value1=32'd15;value2=32'd17;
#400 value1=32'd21;value2=32'd22;
#400 value1=32'd23;value2=32'd26;
#400 value1=32'd37;value2=32'd67;
#400 value1=32'd75;value2=32'd82;
#400 value1=32'd93;value2=32'd116;
#400 value1=32'd217;value2=32'd227;
#400 value1=32'd251;value2=32'd262;
#400 value1=32'd16;value2=32'd18;
#400 value1=32'd21;value2=32'd22;
#400 value1=32'd24;value2=32'd25;
#400 value1=32'd38;value2=32'd68;
#400 value1=32'd76;value2=32'd83;
#400 value1=32'd94;value2=32'd117;
#400 value1=32'd218;value2=32'd228;
#400 value1=32'd252;value2=32'd263;
#400 value1=32'd1;value2=32'd2;
#400 value1=32'd15;value2=32'd28;
#400 value1=32'd29;value2=32'd35;
#400 value1=32'd37;value2=32'd40;
#400 value1=32'd41;value2=32'd43;
#400 value1=32'd45;value2=32'd118;
#400 value1=32'd196;value2=32'd274;
#400 value1=32'd277;value2=32'd279;
#400 value1=32'd1;value2=32'd3;
#400 value1=32'd16;value2=32'd27;
#400 value1=32'd30;value2=32'd36;
#400 value1=32'd38;value2=32'd50;
#400 value1=32'd51;value2=32'd53;
#400 value1=32'd55;value2=32'd119;
#400 value1=32'd197;value2=32'd274;
#400 value1=32'd287;value2=32'd289;
#400 value1=32'd4;value2=32'd14;
#400 value1=32'd17;value2=32'd27;
#400 value1=32'd30;value2=32'd35;
#400 value1=32'd37;value2=32'd60;
#400 value1=32'd62;value2=32'd64;
#400 value1=32'd120;value2=32'd198;
#400 value1=32'd275;value2=32'd285;
#400 value1=32'd296;value2=32'd298;
#400 value1=32'd5;value2=32'd14;
#400 value1=32'd18;value2=32'd28;
#400 value1=32'd29;value2=32'd36;
#400 value1=32'd38;value2=32'd60;
#400 value1=32'd70;value2=32'd72;
#400 value1=32'd121;value2=32'd199;
#400 value1=32'd276;value2=32'd286;
#400 value1=32'd304;value2=32'd306;
#400 value1=32'd6;value2=32'd14;
#400 value1=32'd19;value2=32'd32;
#400 value1=32'd33;value2=32'd35;
#400 value1=32'd36;value2=32'd61;
#400 value1=32'd69;value2=32'd77;
#400 value1=32'd79;value2=32'd122;
#400 value1=32'd200;value2=32'd277;
#400 value1=32'd287;value2=32'd313;
#400 value1=32'd1;value2=32'd7;
#400 value1=32'd20;value2=32'd31;
#400 value1=32'd34;value2=32'd35;
#400 value1=32'd36;value2=32'd62;
#400 value1=32'd70;value2=32'd85;
#400 value1=32'd123;value2=32'd201;
#400 value1=32'd278;value2=32'd288;
#400 value1=32'd312;value2=32'd319;
#400 value1=32'd8;value2=32'd14;
#400 value1=32'd21;value2=32'd31;
#400 value1=32'd34;value2=32'd37;
#400 value1=32'd38;value2=32'd63;
#400 value1=32'd71;value2=32'd84;
#400 value1=32'd90;value2=32'd124;
#400 value1=32'd202;value2=32'd279;
#400 value1=32'd289;value2=32'd313;
#400 value1=32'd1;value2=32'd9;
#400 value1=32'd22;value2=32'd32;
#400 value1=32'd33;value2=32'd37;
#400 value1=32'd38;value2=32'd64;
#400 value1=32'd72;value2=32'd85;
#400 value1=32'd125;value2=32'd203;
#400 value1=32'd280;value2=32'd290;
#400 value1=32'd314;value2=32'd325;
#400 value1=32'd10;value2=32'd23;
#400 value1=32'd27;value2=32'd29;
#400 value1=32'd31;value2=32'd32;
#400 value1=32'd36;value2=32'd37;
#400 value1=32'd65;value2=32'd73;
#400 value1=32'd86;value2=32'd95;
#400 value1=32'd126;value2=32'd204;
#400 value1=32'd281;value2=32'd291;
#400 value1=32'd315;value2=32'd326;
#400 value1=32'd11;value2=32'd24;
#400 value1=32'd28;value2=32'd30;
#400 value1=32'd31;value2=32'd32;
#400 value1=32'd35;value2=32'd38;
#400 value1=32'd66;value2=32'd74;
#400 value1=32'd87;value2=32'd96;
#400 value1=32'd127;value2=32'd205;
#400 value1=32'd282;value2=32'd292;
#400 value1=32'd316;value2=32'd327;
#400 value1=32'd12;value2=32'd25;
#400 value1=32'd27;value2=32'd29;
#400 value1=32'd33;value2=32'd34;
#400 value1=32'd35;value2=32'd38;
#400 value1=32'd67;value2=32'd75;
#400 value1=32'd88;value2=32'd97;
#400 value1=32'd128;value2=32'd206;
#400 value1=32'd283;value2=32'd293;
#400 value1=32'd317;value2=32'd328;
#400 value1=32'd13;value2=32'd26;
#400 value1=32'd28;value2=32'd30;
#400 value1=32'd33;value2=32'd34;
#400 value1=32'd36;value2=32'd37;
#400 value1=32'd68;value2=32'd76;
#400 value1=32'd89;value2=32'd98;
#400 value1=32'd129;value2=32'd207;
#400 value1=32'd284;value2=32'd294;
#400 value1=32'd318;value2=32'd329;
#400 value1=32'd2;value2=32'd3;
#400 value1=32'd41;value2=32'd47;
#400 value1=32'd49;value2=32'd50;
#400 value1=32'd56;value2=32'd58;
#400 value1=32'd130;value2=32'd208;
#400 value1=32'd342;value2=32'd344;
#400 value1=32'd4;value2=32'd15;
#400 value1=32'd27;value2=32'd41;
#400 value1=32'd46;value2=32'd48;
#400 value1=32'd50;value2=32'd65;
#400 value1=32'd67;value2=32'd131;
#400 value1=32'd209;value2=32'd340;
#400 value1=32'd351;value2=32'd353;
#400 value1=32'd5;value2=32'd15;
#400 value1=32'd27;value2=32'd39;
#400 value1=32'd40;value2=32'd47;
#400 value1=32'd49;value2=32'd51;
#400 value1=32'd60;value2=32'd73;
#400 value1=32'd75;value2=32'd132;
#400 value1=32'd210;value2=32'd341;
#400 value1=32'd359;value2=32'd361;
#400 value1=32'd6;value2=32'd15;
#400 value1=32'd43;value2=32'd44;
#400 value1=32'd46;value2=32'd47;
#400 value1=32'd52;value2=32'd61;
#400 value1=32'd80;value2=32'd82;
#400 value1=32'd133;value2=32'd211;
#400 value1=32'd342;value2=32'd368;
#400 value1=32'd2;value2=32'd7;
#400 value1=32'd27;value2=32'd42;
#400 value1=32'd45;value2=32'd46;
#400 value1=32'd47;value2=32'd53;
#400 value1=32'd62;value2=32'd86;
#400 value1=32'd88;value2=32'd134;
#400 value1=32'd212;value2=32'd343;
#400 value1=32'd367;value2=32'd374;
#400 value1=32'd8;value2=32'd15;
#400 value1=32'd42;value2=32'd45;
#400 value1=32'd48;value2=32'd49;
#400 value1=32'd54;value2=32'd63;
#400 value1=32'd91;value2=32'd93;
#400 value1=32'd135;value2=32'd213;
#400 value1=32'd344;value2=32'd368;
#400 value1=32'd2;value2=32'd9;
#400 value1=32'd27;value2=32'd43;
#400 value1=32'd44;value2=32'd48;
#400 value1=32'd49;value2=32'd55;
#400 value1=32'd64;value2=32'd95;
#400 value1=32'd97;value2=32'd136;
#400 value1=32'd214;value2=32'd345;
#400 value1=32'd369;value2=32'd380;
#400 value1=32'd10;value2=32'd40;
#400 value1=32'd42;value2=32'd43;
#400 value1=32'd47;value2=32'd48;
#400 value1=32'd56;value2=32'd65;
#400 value1=32'd100;value2=32'd137;
#400 value1=32'd215;value2=32'd346;
#400 value1=32'd370;value2=32'd381;
#400 value1=32'd11;value2=32'd39;
#400 value1=32'd41;value2=32'd42;
#400 value1=32'd43;value2=32'd46;
#400 value1=32'd49;value2=32'd57;
#400 value1=32'd66;value2=32'd99;
#400 value1=32'd102;value2=32'd138;
#400 value1=32'd216;value2=32'd347;
#400 value1=32'd371;value2=32'd382;
#400 value1=32'd12;value2=32'd40;
#400 value1=32'd44;value2=32'd45;
#400 value1=32'd46;value2=32'd49;
#400 value1=32'd58;value2=32'd67;
#400 value1=32'd100;value2=32'd139;
#400 value1=32'd217;value2=32'd348;
#400 value1=32'd372;value2=32'd383;
#400 value1=32'd13;value2=32'd39;
#400 value1=32'd41;value2=32'd44;
#400 value1=32'd45;value2=32'd47;
#400 value1=32'd48;value2=32'd59;
#400 value1=32'd68;value2=32'd101;
#400 value1=32'd104;value2=32'd140;
#400 value1=32'd218;value2=32'd349;
#400 value1=32'd373;value2=32'd384;
#400 value1=32'd4;value2=32'd16;
#400 value1=32'd28;value2=32'd39;
#400 value1=32'd40;value2=32'd51;
#400 value1=32'd56;value2=32'd58;
#400 value1=32'd60;value2=32'd66;
#400 value1=32'd68;value2=32'd141;
#400 value1=32'd219;value2=32'd340;
#400 value1=32'd396;value2=32'd398;
#400 value1=32'd5;value2=32'd16;
#400 value1=32'd28;value2=32'd41;
#400 value1=32'd50;value2=32'd57;
#400 value1=32'd59;value2=32'd74;
#400 value1=32'd76;value2=32'd142;
#400 value1=32'd220;value2=32'd341;
#400 value1=32'd404;value2=32'd406;
#400 value1=32'd6;value2=32'd16;
#400 value1=32'd42;value2=32'd53;
#400 value1=32'd54;value2=32'd56;
#400 value1=32'd57;value2=32'd69;
#400 value1=32'd81;value2=32'd83;
#400 value1=32'd143;value2=32'd221;
#400 value1=32'd342;value2=32'd413;
#400 value1=32'd3;value2=32'd7;
#400 value1=32'd28;value2=32'd43;
#400 value1=32'd52;value2=32'd55;
#400 value1=32'd56;value2=32'd57;
#400 value1=32'd70;value2=32'd87;
#400 value1=32'd89;value2=32'd144;
#400 value1=32'd222;value2=32'd343;
#400 value1=32'd412;value2=32'd419;
#400 value1=32'd8;value2=32'd16;
#400 value1=32'd44;value2=32'd52;
#400 value1=32'd55;value2=32'd58;
#400 value1=32'd59;value2=32'd71;
#400 value1=32'd92;value2=32'd94;
#400 value1=32'd145;value2=32'd223;
#400 value1=32'd344;value2=32'd413;
#400 value1=32'd3;value2=32'd9;
#400 value1=32'd28;value2=32'd45;
#400 value1=32'd53;value2=32'd54;
#400 value1=32'd58;value2=32'd59;
#400 value1=32'd72;value2=32'd96;
#400 value1=32'd98;value2=32'd146;
#400 value1=32'd224;value2=32'd345;
#400 value1=32'd414;value2=32'd425;
#400 value1=32'd10;value2=32'd39;
#400 value1=32'd46;value2=32'd50;
#400 value1=32'd52;value2=32'd53;
#400 value1=32'd57;value2=32'd58;
#400 value1=32'd73;value2=32'd99;
#400 value1=32'd101;value2=32'd147;
#400 value1=32'd225;value2=32'd346;
#400 value1=32'd415;value2=32'd426;
#400 value1=32'd11;value2=32'd47;
#400 value1=32'd51;value2=32'd52;
#400 value1=32'd53;value2=32'd56;
#400 value1=32'd59;value2=32'd74;
#400 value1=32'd103;value2=32'd148;
#400 value1=32'd226;value2=32'd347;
#400 value1=32'd416;value2=32'd427;
#400 value1=32'd12;value2=32'd39;
#400 value1=32'd48;value2=32'd50;
#400 value1=32'd54;value2=32'd55;
#400 value1=32'd56;value2=32'd59;
#400 value1=32'd75;value2=32'd102;
#400 value1=32'd104;value2=32'd149;
#400 value1=32'd227;value2=32'd348;
#400 value1=32'd417;value2=32'd428;
#400 value1=32'd13;value2=32'd49;
#400 value1=32'd51;value2=32'd54;
#400 value1=32'd55;value2=32'd57;
#400 value1=32'd58;value2=32'd76;
#400 value1=32'd103;value2=32'd150;
#400 value1=32'd228;value2=32'd349;
#400 value1=32'd418;value2=32'd429;
#400 value1=32'd17;value2=32'd18;
#400 value1=32'd29;value2=32'd30;
#400 value1=32'd41;value2=32'd50;
#400 value1=32'd66;value2=32'd68;
#400 value1=32'd73;value2=32'd75;
#400 value1=32'd151;value2=32'd229;
#400 value1=32'd350;value2=32'd395;
#400 value1=32'd440;value2=32'd442;
#400 value1=32'd17;value2=32'd19;
#400 value1=32'd31;value2=32'd42;
#400 value1=32'd62;value2=32'd63;
#400 value1=32'd65;value2=32'd66;
#400 value1=32'd69;value2=32'd80;
#400 value1=32'd82;value2=32'd152;
#400 value1=32'd230;value2=32'd351;
#400 value1=32'd396;value2=32'd449;
#400 value1=32'd4;value2=32'd20;
#400 value1=32'd29;value2=32'd32;
#400 value1=32'd43;value2=32'd61;
#400 value1=32'd64;value2=32'd65;
#400 value1=32'd66;value2=32'd70;
#400 value1=32'd86;value2=32'd88;
#400 value1=32'd153;value2=32'd231;
#400 value1=32'd352;value2=32'd397;
#400 value1=32'd448;value2=32'd455;
#400 value1=32'd17;value2=32'd21;
#400 value1=32'd33;value2=32'd44;
#400 value1=32'd61;value2=32'd64;
#400 value1=32'd67;value2=32'd68;
#400 value1=32'd71;value2=32'd91;
#400 value1=32'd93;value2=32'd154;
#400 value1=32'd232;value2=32'd353;
#400 value1=32'd398;value2=32'd449;
#400 value1=32'd4;value2=32'd22;
#400 value1=32'd29;value2=32'd34;
#400 value1=32'd45;value2=32'd62;
#400 value1=32'd63;value2=32'd67;
#400 value1=32'd68;value2=32'd72;
#400 value1=32'd95;value2=32'd97;
#400 value1=32'd155;value2=32'd233;
#400 value1=32'd354;value2=32'd399;
#400 value1=32'd450;value2=32'd461;
#400 value1=32'd23;value2=32'd35;
#400 value1=32'd40;value2=32'd46;
#400 value1=32'd61;value2=32'd62;
#400 value1=32'd66;value2=32'd67;
#400 value1=32'd73;value2=32'd100;
#400 value1=32'd156;value2=32'd234;
#400 value1=32'd355;value2=32'd400;
#400 value1=32'd451;value2=32'd462;
#400 value1=32'd24;value2=32'd36;
#400 value1=32'd47;value2=32'd50;
#400 value1=32'd60;value2=32'd61;
#400 value1=32'd62;value2=32'd65;
#400 value1=32'd68;value2=32'd74;
#400 value1=32'd99;value2=32'd102;
#400 value1=32'd157;value2=32'd235;
#400 value1=32'd356;value2=32'd401;
#400 value1=32'd452;value2=32'd463;
#400 value1=32'd25;value2=32'd37;
#400 value1=32'd40;value2=32'd48;
#400 value1=32'd63;value2=32'd64;
#400 value1=32'd65;value2=32'd68;
#400 value1=32'd75;value2=32'd100;
#400 value1=32'd158;value2=32'd236;
#400 value1=32'd357;value2=32'd402;
#400 value1=32'd453;value2=32'd464;
#400 value1=32'd26;value2=32'd38;
#400 value1=32'd49;value2=32'd50;
#400 value1=32'd60;value2=32'd63;
#400 value1=32'd64;value2=32'd66;
#400 value1=32'd67;value2=32'd76;
#400 value1=32'd101;value2=32'd104;
#400 value1=32'd159;value2=32'd237;
#400 value1=32'd358;value2=32'd403;
#400 value1=32'd454;value2=32'd465;
#400 value1=32'd18;value2=32'd19;
#400 value1=32'd31;value2=32'd52;
#400 value1=32'd61;value2=32'd70;
#400 value1=32'd71;value2=32'd73;
#400 value1=32'd74;value2=32'd81;
#400 value1=32'd83;value2=32'd160;
#400 value1=32'd238;value2=32'd359;
#400 value1=32'd404;value2=32'd477;
#400 value1=32'd5;value2=32'd20;
#400 value1=32'd30;value2=32'd32;
#400 value1=32'd53;value2=32'd62;
#400 value1=32'd69;value2=32'd72;
#400 value1=32'd73;value2=32'd74;
#400 value1=32'd87;value2=32'd89;
#400 value1=32'd161;value2=32'd239;
#400 value1=32'd360;value2=32'd405;
#400 value1=32'd476;value2=32'd483;
#400 value1=32'd18;value2=32'd21;
#400 value1=32'd33;value2=32'd54;
#400 value1=32'd63;value2=32'd69;
#400 value1=32'd72;value2=32'd75;
#400 value1=32'd76;value2=32'd92;
#400 value1=32'd94;value2=32'd162;
#400 value1=32'd240;value2=32'd361;
#400 value1=32'd406;value2=32'd477;
#400 value1=32'd5;value2=32'd22;
#400 value1=32'd30;value2=32'd34;
#400 value1=32'd55;value2=32'd64;
#400 value1=32'd70;value2=32'd71;
#400 value1=32'd75;value2=32'd76;
#400 value1=32'd96;value2=32'd98;
#400 value1=32'd163;value2=32'd241;
#400 value1=32'd362;value2=32'd407;
#400 value1=32'd478;value2=32'd489;
#400 value1=32'd23;value2=32'd35;
#400 value1=32'd41;value2=32'd56;
#400 value1=32'd60;value2=32'd65;
#400 value1=32'd69;value2=32'd70;
#400 value1=32'd74;value2=32'd75;
#400 value1=32'd99;value2=32'd101;
#400 value1=32'd164;value2=32'd242;
#400 value1=32'd363;value2=32'd408;
#400 value1=32'd479;value2=32'd490;
#400 value1=32'd24;value2=32'd36;
#400 value1=32'd51;value2=32'd57;
#400 value1=32'd66;value2=32'd69;
#400 value1=32'd70;value2=32'd73;
#400 value1=32'd76;value2=32'd103;
#400 value1=32'd165;value2=32'd243;
#400 value1=32'd364;value2=32'd409;
#400 value1=32'd480;value2=32'd491;
#400 value1=32'd25;value2=32'd37;
#400 value1=32'd41;value2=32'd58;
#400 value1=32'd60;value2=32'd67;
#400 value1=32'd71;value2=32'd72;
#400 value1=32'd73;value2=32'd76;
#400 value1=32'd102;value2=32'd104;
#400 value1=32'd166;value2=32'd244;
#400 value1=32'd365;value2=32'd410;
#400 value1=32'd481;value2=32'd492;
#400 value1=32'd26;value2=32'd38;
#400 value1=32'd51;value2=32'd59;
#400 value1=32'd68;value2=32'd71;
#400 value1=32'd72;value2=32'd74;
#400 value1=32'd75;value2=32'd103;
#400 value1=32'd167;value2=32'd245;
#400 value1=32'd366;value2=32'd411;
#400 value1=32'd482;value2=32'd493;
#400 value1=32'd6;value2=32'd20;
#400 value1=32'd31;value2=32'd79;
#400 value1=32'd80;value2=32'd81;
#400 value1=32'd84;value2=32'd86;
#400 value1=32'd87;value2=32'd168;
#400 value1=32'd246;value2=32'd367;
#400 value1=32'd412;value2=32'd504;
#400 value1=32'd19;value2=32'd21;
#400 value1=32'd79;value2=32'd82;
#400 value1=32'd83;value2=32'd84;
#400 value1=32'd91;value2=32'd92;
#400 value1=32'd169;value2=32'd247;
#400 value1=32'd368;value2=32'd413;
#400 value1=32'd6;value2=32'd22;
#400 value1=32'd31;value2=32'd77;
#400 value1=32'd78;value2=32'd82;
#400 value1=32'd83;value2=32'd85;
#400 value1=32'd90;value2=32'd95;
#400 value1=32'd96;value2=32'd170;
#400 value1=32'd248;value2=32'd369;
#400 value1=32'd414;value2=32'd510;
#400 value1=32'd23;value2=32'd42;
#400 value1=32'd61;value2=32'd77;
#400 value1=32'd81;value2=32'd82;
#400 value1=32'd86;value2=32'd91;
#400 value1=32'd99;value2=32'd171;
#400 value1=32'd249;value2=32'd370;
#400 value1=32'd415;value2=32'd511;
#400 value1=32'd24;value2=32'd52;
#400 value1=32'd69;value2=32'd77;
#400 value1=32'd80;value2=32'd83;
#400 value1=32'd87;value2=32'd92;
#400 value1=32'd99;value2=32'd172;
#400 value1=32'd250;value2=32'd371;
#400 value1=32'd416;value2=32'd512;
#400 value1=32'd25;value2=32'd42;
#400 value1=32'd61;value2=32'd78;
#400 value1=32'd79;value2=32'd80;
#400 value1=32'd83;value2=32'd88;
#400 value1=32'd93;value2=32'd100;
#400 value1=32'd102;value2=32'd173;
#400 value1=32'd251;value2=32'd372;
#400 value1=32'd417;value2=32'd513;
#400 value1=32'd26;value2=32'd52;
#400 value1=32'd69;value2=32'd78;
#400 value1=32'd79;value2=32'd81;
#400 value1=32'd82;value2=32'd89;
#400 value1=32'd94;value2=32'd101;
#400 value1=32'd103;value2=32'd174;
#400 value1=32'd252;value2=32'd373;
#400 value1=32'd418;value2=32'd514;
#400 value1=32'd8;value2=32'd20;
#400 value1=32'd33;value2=32'd77;
#400 value1=32'd78;value2=32'd85;
#400 value1=32'd88;value2=32'd89;
#400 value1=32'd90;value2=32'd91;
#400 value1=32'd92;value2=32'd175;
#400 value1=32'd253;value2=32'd374;
#400 value1=32'd419;value2=32'd504;
#400 value1=32'd7;value2=32'd9;
#400 value1=32'd32;value2=32'd34;
#400 value1=32'd79;value2=32'd84;
#400 value1=32'd88;value2=32'd89;
#400 value1=32'd95;value2=32'd96;
#400 value1=32'd176;value2=32'd254;
#400 value1=32'd375;value2=32'd420;
#400 value1=32'd505;value2=32'd525;
#400 value1=32'd10;value2=32'd35;
#400 value1=32'd43;value2=32'd62;
#400 value1=32'd77;value2=32'd80;
#400 value1=32'd87;value2=32'd88;
#400 value1=32'd95;value2=32'd99;
#400 value1=32'd177;value2=32'd255;
#400 value1=32'd376;value2=32'd421;
#400 value1=32'd506;value2=32'd526;
#400 value1=32'd11;value2=32'd36;
#400 value1=32'd53;value2=32'd70;
#400 value1=32'd77;value2=32'd81;
#400 value1=32'd86;value2=32'd89;
#400 value1=32'd96;value2=32'd99;
#400 value1=32'd178;value2=32'd256;
#400 value1=32'd377;value2=32'd422;
#400 value1=32'd507;value2=32'd527;
#400 value1=32'd12;value2=32'd37;
#400 value1=32'd43;value2=32'd62;
#400 value1=32'd82;value2=32'd84;
#400 value1=32'd85;value2=32'd86;
#400 value1=32'd89;value2=32'd97;
#400 value1=32'd100;value2=32'd102;
#400 value1=32'd179;value2=32'd257;
#400 value1=32'd378;value2=32'd423;
#400 value1=32'd508;value2=32'd528;
#400 value1=32'd13;value2=32'd38;
#400 value1=32'd53;value2=32'd70;
#400 value1=32'd83;value2=32'd84;
#400 value1=32'd85;value2=32'd87;
#400 value1=32'd88;value2=32'd98;
#400 value1=32'd101;value2=32'd103;
#400 value1=32'd180;value2=32'd258;
#400 value1=32'd379;value2=32'd424;
#400 value1=32'd509;value2=32'd529;
#400 value1=32'd8;value2=32'd22;
#400 value1=32'd33;value2=32'd79;
#400 value1=32'd84;value2=32'd93;
#400 value1=32'd94;value2=32'd97;
#400 value1=32'd98;value2=32'd181;
#400 value1=32'd259;value2=32'd380;
#400 value1=32'd425;value2=32'd510;
#400 value1=32'd23;value2=32'd44;
#400 value1=32'd63;value2=32'd78;
#400 value1=32'd80;value2=32'd84;
#400 value1=32'd92;value2=32'd93;
#400 value1=32'd95;value2=32'd100;
#400 value1=32'd101;value2=32'd182;
#400 value1=32'd260;value2=32'd381;
#400 value1=32'd426;value2=32'd511;
#400 value1=32'd24;value2=32'd54;
#400 value1=32'd71;value2=32'd78;
#400 value1=32'd81;value2=32'd84;
#400 value1=32'd91;value2=32'd94;
#400 value1=32'd96;value2=32'd102;
#400 value1=32'd103;value2=32'd183;
#400 value1=32'd261;value2=32'd382;
#400 value1=32'd427;value2=32'd512;
#400 value1=32'd25;value2=32'd44;
#400 value1=32'd63;value2=32'd82;
#400 value1=32'd90;value2=32'd91;
#400 value1=32'd94;value2=32'd97;
#400 value1=32'd104;value2=32'd184;
#400 value1=32'd262;value2=32'd383;
#400 value1=32'd428;value2=32'd513;
#400 value1=32'd26;value2=32'd54;
#400 value1=32'd71;value2=32'd83;
#400 value1=32'd90;value2=32'd92;
#400 value1=32'd93;value2=32'd98;
#400 value1=32'd104;value2=32'd185;
#400 value1=32'd263;value2=32'd384;
#400 value1=32'd429;value2=32'd514;
#400 value1=32'd10;value2=32'd35;
#400 value1=32'd45;value2=32'd64;
#400 value1=32'd79;value2=32'd85;
#400 value1=32'd86;value2=32'd91;
#400 value1=32'd96;value2=32'd97;
#400 value1=32'd100;value2=32'd101;
#400 value1=32'd186;value2=32'd264;
#400 value1=32'd385;value2=32'd430;
#400 value1=32'd515;value2=32'd540;
#400 value1=32'd11;value2=32'd36;
#400 value1=32'd55;value2=32'd72;
#400 value1=32'd79;value2=32'd85;
#400 value1=32'd87;value2=32'd92;
#400 value1=32'd95;value2=32'd98;
#400 value1=32'd102;value2=32'd103;
#400 value1=32'd187;value2=32'd265;
#400 value1=32'd386;value2=32'd431;
#400 value1=32'd516;value2=32'd541;
#400 value1=32'd12;value2=32'd37;
#400 value1=32'd45;value2=32'd64;
#400 value1=32'd88;value2=32'd90;
#400 value1=32'd93;value2=32'd95;
#400 value1=32'd98;value2=32'd104;
#400 value1=32'd188;value2=32'd266;
#400 value1=32'd387;value2=32'd432;
#400 value1=32'd517;value2=32'd542;
#400 value1=32'd13;value2=32'd38;
#400 value1=32'd55;value2=32'd72;
#400 value1=32'd89;value2=32'd90;
#400 value1=32'd94;value2=32'd96;
#400 value1=32'd97;value2=32'd104;
#400 value1=32'd189;value2=32'd267;
#400 value1=32'd388;value2=32'd433;
#400 value1=32'd518;value2=32'd543;
#400 value1=32'd47;value2=32'd56;
#400 value1=32'd66;value2=32'd73;
#400 value1=32'd80;value2=32'd81;
#400 value1=32'd86;value2=32'd87;
#400 value1=32'd101;value2=32'd102;
#400 value1=32'd190;value2=32'd268;
#400 value1=32'd389;value2=32'd434;
#400 value1=32'd519;value2=32'd544;
#400 value1=32'd46;value2=32'd48;
#400 value1=32'd65;value2=32'd67;
#400 value1=32'd82;value2=32'd88;
#400 value1=32'd91;value2=32'd95;
#400 value1=32'd101;value2=32'd102;
#400 value1=32'd191;value2=32'd269;
#400 value1=32'd390;value2=32'd435;
#400 value1=32'd520;value2=32'd545;
#400 value1=32'd49;value2=32'd56;
#400 value1=32'd68;value2=32'd73;
#400 value1=32'd83;value2=32'd89;
#400 value1=32'd91;value2=32'd95;
#400 value1=32'd99;value2=32'd100;
#400 value1=32'd103;value2=32'd104;
#400 value1=32'd192;value2=32'd270;
#400 value1=32'd391;value2=32'd436;
#400 value1=32'd521;value2=32'd546;
#400 value1=32'd47;value2=32'd58;
#400 value1=32'd66;value2=32'd75;
#400 value1=32'd82;value2=32'd88;
#400 value1=32'd92;value2=32'd96;
#400 value1=32'd99;value2=32'd100;
#400 value1=32'd103;value2=32'd104;
#400 value1=32'd193;value2=32'd271;
#400 value1=32'd392;value2=32'd437;
#400 value1=32'd522;value2=32'd547;
#400 value1=32'd57;value2=32'd59;
#400 value1=32'd74;value2=32'd76;
#400 value1=32'd83;value2=32'd89;
#400 value1=32'd92;value2=32'd96;
#400 value1=32'd101;value2=32'd102;
#400 value1=32'd194;value2=32'd272;
#400 value1=32'd393;value2=32'd438;
#400 value1=32'd523;value2=32'd548;
#400 value1=32'd49;value2=32'd58;
#400 value1=32'd68;value2=32'd75;
#400 value1=32'd93;value2=32'd94;
#400 value1=32'd97;value2=32'd98;
#400 value1=32'd101;value2=32'd102;
#400 value1=32'd195;value2=32'd273;
#400 value1=32'd394;value2=32'd439;
#400 value1=32'd524;value2=32'd549;
#400 value1=32'd1;value2=32'd14;
#400 value1=32'd108;value2=32'd109;
#400 value1=32'd111;value2=32'd113;
#400 value1=32'd120;value2=32'd121;
#400 value1=32'd122;value2=32'd124;
#400 value1=32'd196;value2=32'd197;
#400 value1=32'd201;value2=32'd203;
#400 value1=32'd0;value2=32'd2;
#400 value1=32'd15;value2=32'd107;
#400 value1=32'd108;value2=32'd114;
#400 value1=32'd116;value2=32'd118;
#400 value1=32'd131;value2=32'd132;
#400 value1=32'd133;value2=32'd135;
#400 value1=32'd196;value2=32'd208;
#400 value1=32'd212;value2=32'd214;
#400 value1=32'd0;value2=32'd3;
#400 value1=32'd16;value2=32'd106;
#400 value1=32'd109;value2=32'd115;
#400 value1=32'd117;value2=32'd119;
#400 value1=32'd141;value2=32'd142;
#400 value1=32'd143;value2=32'd145;
#400 value1=32'd197;value2=32'd208;
#400 value1=32'd222;value2=32'd224;
#400 value1=32'd4;value2=32'd17;
#400 value1=32'd105;value2=32'd106;
#400 value1=32'd109;value2=32'd114;
#400 value1=32'd116;value2=32'd120;
#400 value1=32'd151;value2=32'd152;
#400 value1=32'd154;value2=32'd198;
#400 value1=32'd209;value2=32'd219;
#400 value1=32'd231;value2=32'd233;
#400 value1=32'd5;value2=32'd18;
#400 value1=32'd105;value2=32'd107;
#400 value1=32'd108;value2=32'd115;
#400 value1=32'd117;value2=32'd121;
#400 value1=32'd151;value2=32'd160;
#400 value1=32'd162;value2=32'd199;
#400 value1=32'd210;value2=32'd220;
#400 value1=32'd239;value2=32'd241;
#400 value1=32'd0;value2=32'd6;
#400 value1=32'd19;value2=32'd111;
#400 value1=32'd112;value2=32'd114;
#400 value1=32'd115;value2=32'd122;
#400 value1=32'd152;value2=32'd160;
#400 value1=32'd169;value2=32'd200;
#400 value1=32'd211;value2=32'd221;
#400 value1=32'd246;value2=32'd248;
#400 value1=32'd7;value2=32'd20;
#400 value1=32'd105;value2=32'd110;
#400 value1=32'd113;value2=32'd114;
#400 value1=32'd115;value2=32'd123;
#400 value1=32'd153;value2=32'd161;
#400 value1=32'd168;value2=32'd175;
#400 value1=32'd201;value2=32'd212;
#400 value1=32'd222;value2=32'd254;
#400 value1=32'd0;value2=32'd8;
#400 value1=32'd21;value2=32'd110;
#400 value1=32'd113;value2=32'd116;
#400 value1=32'd117;value2=32'd124;
#400 value1=32'd154;value2=32'd162;
#400 value1=32'd169;value2=32'd202;
#400 value1=32'd213;value2=32'd223;
#400 value1=32'd253;value2=32'd259;
#400 value1=32'd9;value2=32'd22;
#400 value1=32'd105;value2=32'd111;
#400 value1=32'd112;value2=32'd116;
#400 value1=32'd117;value2=32'd125;
#400 value1=32'd155;value2=32'd163;
#400 value1=32'd170;value2=32'd181;
#400 value1=32'd203;value2=32'd214;
#400 value1=32'd224;value2=32'd254;
#400 value1=32'd10;value2=32'd23;
#400 value1=32'd106;value2=32'd108;
#400 value1=32'd110;value2=32'd111;
#400 value1=32'd115;value2=32'd116;
#400 value1=32'd126;value2=32'd156;
#400 value1=32'd164;value2=32'd171;
#400 value1=32'd182;value2=32'd204;
#400 value1=32'd215;value2=32'd225;
#400 value1=32'd255;value2=32'd264;
#400 value1=32'd11;value2=32'd24;
#400 value1=32'd107;value2=32'd109;
#400 value1=32'd110;value2=32'd111;
#400 value1=32'd114;value2=32'd117;
#400 value1=32'd127;value2=32'd157;
#400 value1=32'd165;value2=32'd172;
#400 value1=32'd183;value2=32'd205;
#400 value1=32'd216;value2=32'd226;
#400 value1=32'd256;value2=32'd265;
#400 value1=32'd12;value2=32'd25;
#400 value1=32'd106;value2=32'd108;
#400 value1=32'd112;value2=32'd113;
#400 value1=32'd114;value2=32'd117;
#400 value1=32'd128;value2=32'd158;
#400 value1=32'd166;value2=32'd173;
#400 value1=32'd184;value2=32'd206;
#400 value1=32'd217;value2=32'd227;
#400 value1=32'd257;value2=32'd266;
#400 value1=32'd13;value2=32'd26;
#400 value1=32'd107;value2=32'd109;
#400 value1=32'd112;value2=32'd113;
#400 value1=32'd115;value2=32'd116;
#400 value1=32'd129;value2=32'd159;
#400 value1=32'd167;value2=32'd174;
#400 value1=32'd185;value2=32'd207;
#400 value1=32'd218;value2=32'd228;
#400 value1=32'd258;value2=32'd267;
#400 value1=32'd1;value2=32'd27;
#400 value1=32'd106;value2=32'd119;
#400 value1=32'd120;value2=32'd126;
#400 value1=32'd128;value2=32'd131;
#400 value1=32'd132;value2=32'd134;
#400 value1=32'd136;value2=32'd274;
#400 value1=32'd278;value2=32'd280;
#400 value1=32'd1;value2=32'd28;
#400 value1=32'd107;value2=32'd118;
#400 value1=32'd121;value2=32'd127;
#400 value1=32'd129;value2=32'd141;
#400 value1=32'd142;value2=32'd144;
#400 value1=32'd146;value2=32'd274;
#400 value1=32'd288;value2=32'd290;
#400 value1=32'd29;value2=32'd105;
#400 value1=32'd108;value2=32'd118;
#400 value1=32'd121;value2=32'd126;
#400 value1=32'd128;value2=32'd151;
#400 value1=32'd153;value2=32'd155;
#400 value1=32'd275;value2=32'd285;
#400 value1=32'd297;value2=32'd299;
#400 value1=32'd30;value2=32'd105;
#400 value1=32'd109;value2=32'd119;
#400 value1=32'd120;value2=32'd127;
#400 value1=32'd129;value2=32'd151;
#400 value1=32'd161;value2=32'd163;
#400 value1=32'd276;value2=32'd286;
#400 value1=32'd305;value2=32'd307;
#400 value1=32'd1;value2=32'd31;
#400 value1=32'd105;value2=32'd110;
#400 value1=32'd123;value2=32'd124;
#400 value1=32'd126;value2=32'd127;
#400 value1=32'd152;value2=32'd160;
#400 value1=32'd168;value2=32'd170;
#400 value1=32'd277;value2=32'd287;
#400 value1=32'd312;value2=32'd314;
#400 value1=32'd32;value2=32'd111;
#400 value1=32'd122;value2=32'd125;
#400 value1=32'd126;value2=32'd127;
#400 value1=32'd153;value2=32'd161;
#400 value1=32'd176;value2=32'd278;
#400 value1=32'd288;value2=32'd320;
#400 value1=32'd1;value2=32'd33;
#400 value1=32'd105;value2=32'd112;
#400 value1=32'd122;value2=32'd125;
#400 value1=32'd128;value2=32'd129;
#400 value1=32'd154;value2=32'd162;
#400 value1=32'd175;value2=32'd181;
#400 value1=32'd279;value2=32'd289;
#400 value1=32'd319;value2=32'd325;
#400 value1=32'd34;value2=32'd113;
#400 value1=32'd123;value2=32'd124;
#400 value1=32'd128;value2=32'd129;
#400 value1=32'd155;value2=32'd163;
#400 value1=32'd176;value2=32'd280;
#400 value1=32'd290;value2=32'd320;
#400 value1=32'd35;value2=32'd114;
#400 value1=32'd118;value2=32'd120;
#400 value1=32'd122;value2=32'd123;
#400 value1=32'd127;value2=32'd128;
#400 value1=32'd156;value2=32'd164;
#400 value1=32'd177;value2=32'd186;
#400 value1=32'd281;value2=32'd291;
#400 value1=32'd321;value2=32'd330;
#400 value1=32'd36;value2=32'd115;
#400 value1=32'd119;value2=32'd121;
#400 value1=32'd122;value2=32'd123;
#400 value1=32'd126;value2=32'd129;
#400 value1=32'd157;value2=32'd165;
#400 value1=32'd178;value2=32'd187;
#400 value1=32'd282;value2=32'd292;
#400 value1=32'd322;value2=32'd331;
#400 value1=32'd37;value2=32'd116;
#400 value1=32'd118;value2=32'd120;
#400 value1=32'd124;value2=32'd125;
#400 value1=32'd126;value2=32'd129;
#400 value1=32'd158;value2=32'd166;
#400 value1=32'd179;value2=32'd188;
#400 value1=32'd283;value2=32'd293;
#400 value1=32'd323;value2=32'd332;
#400 value1=32'd38;value2=32'd117;
#400 value1=32'd119;value2=32'd121;
#400 value1=32'd124;value2=32'd125;
#400 value1=32'd127;value2=32'd128;
#400 value1=32'd159;value2=32'd167;
#400 value1=32'd180;value2=32'd189;
#400 value1=32'd284;value2=32'd294;
#400 value1=32'd324;value2=32'd333;
#400 value1=32'd2;value2=32'd3;
#400 value1=32'd39;value2=32'd132;
#400 value1=32'd138;value2=32'd140;
#400 value1=32'd141;value2=32'd147;
#400 value1=32'd149;value2=32'd274;
#400 value1=32'd343;value2=32'd345;
#400 value1=32'd4;value2=32'd40;
#400 value1=32'd106;value2=32'd118;
#400 value1=32'd132;value2=32'd137;
#400 value1=32'd139;value2=32'd141;
#400 value1=32'd156;value2=32'd158;
#400 value1=32'd275;value2=32'd340;
#400 value1=32'd352;value2=32'd354;
#400 value1=32'd5;value2=32'd41;
#400 value1=32'd106;value2=32'd118;
#400 value1=32'd130;value2=32'd131;
#400 value1=32'd138;value2=32'd140;
#400 value1=32'd142;value2=32'd151;
#400 value1=32'd164;value2=32'd166;
#400 value1=32'd276;value2=32'd341;
#400 value1=32'd360;value2=32'd362;
#400 value1=32'd2;value2=32'd6;
#400 value1=32'd42;value2=32'd106;
#400 value1=32'd134;value2=32'd135;
#400 value1=32'd137;value2=32'd138;
#400 value1=32'd143;value2=32'd152;
#400 value1=32'd171;value2=32'd173;
#400 value1=32'd277;value2=32'd342;
#400 value1=32'd367;value2=32'd369;
#400 value1=32'd7;value2=32'd43;
#400 value1=32'd118;value2=32'd133;
#400 value1=32'd136;value2=32'd137;
#400 value1=32'd138;value2=32'd144;
#400 value1=32'd153;value2=32'd177;
#400 value1=32'd179;value2=32'd278;
#400 value1=32'd343;value2=32'd375;
#400 value1=32'd2;value2=32'd8;
#400 value1=32'd44;value2=32'd106;
#400 value1=32'd133;value2=32'd136;
#400 value1=32'd139;value2=32'd140;
#400 value1=32'd145;value2=32'd154;
#400 value1=32'd182;value2=32'd184;
#400 value1=32'd279;value2=32'd344;
#400 value1=32'd374;value2=32'd380;
#400 value1=32'd9;value2=32'd45;
#400 value1=32'd118;value2=32'd134;
#400 value1=32'd135;value2=32'd139;
#400 value1=32'd140;value2=32'd146;
#400 value1=32'd155;value2=32'd186;
#400 value1=32'd188;value2=32'd280;
#400 value1=32'd345;value2=32'd375;
#400 value1=32'd10;value2=32'd46;
#400 value1=32'd131;value2=32'd133;
#400 value1=32'd134;value2=32'd138;
#400 value1=32'd139;value2=32'd147;
#400 value1=32'd156;value2=32'd191;
#400 value1=32'd281;value2=32'd346;
#400 value1=32'd376;value2=32'd385;
#400 value1=32'd11;value2=32'd47;
#400 value1=32'd130;value2=32'd132;
#400 value1=32'd133;value2=32'd134;
#400 value1=32'd137;value2=32'd140;
#400 value1=32'd148;value2=32'd157;
#400 value1=32'd190;value2=32'd193;
#400 value1=32'd282;value2=32'd347;
#400 value1=32'd377;value2=32'd386;
#400 value1=32'd12;value2=32'd48;
#400 value1=32'd131;value2=32'd135;
#400 value1=32'd136;value2=32'd137;
#400 value1=32'd140;value2=32'd149;
#400 value1=32'd158;value2=32'd191;
#400 value1=32'd283;value2=32'd348;
#400 value1=32'd378;value2=32'd387;
#400 value1=32'd13;value2=32'd49;
#400 value1=32'd130;value2=32'd132;
#400 value1=32'd135;value2=32'd136;
#400 value1=32'd138;value2=32'd139;
#400 value1=32'd150;value2=32'd159;
#400 value1=32'd192;value2=32'd195;
#400 value1=32'd284;value2=32'd349;
#400 value1=32'd379;value2=32'd388;
#400 value1=32'd4;value2=32'd50;
#400 value1=32'd107;value2=32'd119;
#400 value1=32'd130;value2=32'd131;
#400 value1=32'd142;value2=32'd147;
#400 value1=32'd149;value2=32'd151;
#400 value1=32'd157;value2=32'd159;
#400 value1=32'd285;value2=32'd340;
#400 value1=32'd397;value2=32'd399;
#400 value1=32'd5;value2=32'd51;
#400 value1=32'd107;value2=32'd119;
#400 value1=32'd132;value2=32'd141;
#400 value1=32'd148;value2=32'd150;
#400 value1=32'd165;value2=32'd167;
#400 value1=32'd286;value2=32'd341;
#400 value1=32'd405;value2=32'd407;
#400 value1=32'd3;value2=32'd6;
#400 value1=32'd52;value2=32'd107;
#400 value1=32'd133;value2=32'd144;
#400 value1=32'd145;value2=32'd147;
#400 value1=32'd148;value2=32'd160;
#400 value1=32'd172;value2=32'd174;
#400 value1=32'd287;value2=32'd342;
#400 value1=32'd412;value2=32'd414;
#400 value1=32'd7;value2=32'd53;
#400 value1=32'd119;value2=32'd134;
#400 value1=32'd143;value2=32'd146;
#400 value1=32'd147;value2=32'd148;
#400 value1=32'd161;value2=32'd178;
#400 value1=32'd180;value2=32'd288;
#400 value1=32'd343;value2=32'd420;
#400 value1=32'd3;value2=32'd8;
#400 value1=32'd54;value2=32'd107;
#400 value1=32'd135;value2=32'd143;
#400 value1=32'd146;value2=32'd149;
#400 value1=32'd150;value2=32'd162;
#400 value1=32'd183;value2=32'd185;
#400 value1=32'd289;value2=32'd344;
#400 value1=32'd419;value2=32'd425;
#400 value1=32'd9;value2=32'd55;
#400 value1=32'd119;value2=32'd136;
#400 value1=32'd144;value2=32'd145;
#400 value1=32'd149;value2=32'd150;
#400 value1=32'd163;value2=32'd187;
#400 value1=32'd189;value2=32'd290;
#400 value1=32'd345;value2=32'd420;
#400 value1=32'd10;value2=32'd56;
#400 value1=32'd130;value2=32'd137;
#400 value1=32'd141;value2=32'd143;
#400 value1=32'd144;value2=32'd148;
#400 value1=32'd149;value2=32'd164;
#400 value1=32'd190;value2=32'd192;
#400 value1=32'd291;value2=32'd346;
#400 value1=32'd421;value2=32'd430;
#400 value1=32'd11;value2=32'd57;
#400 value1=32'd138;value2=32'd142;
#400 value1=32'd143;value2=32'd144;
#400 value1=32'd147;value2=32'd150;
#400 value1=32'd165;value2=32'd194;
#400 value1=32'd292;value2=32'd347;
#400 value1=32'd422;value2=32'd431;
#400 value1=32'd12;value2=32'd58;
#400 value1=32'd130;value2=32'd139;
#400 value1=32'd141;value2=32'd145;
#400 value1=32'd146;value2=32'd147;
#400 value1=32'd150;value2=32'd166;
#400 value1=32'd193;value2=32'd195;
#400 value1=32'd293;value2=32'd348;
#400 value1=32'd423;value2=32'd432;
#400 value1=32'd13;value2=32'd59;
#400 value1=32'd140;value2=32'd142;
#400 value1=32'd145;value2=32'd146;
#400 value1=32'd148;value2=32'd149;
#400 value1=32'd167;value2=32'd194;
#400 value1=32'd294;value2=32'd349;
#400 value1=32'd424;value2=32'd433;
#400 value1=32'd60;value2=32'd108;
#400 value1=32'd109;value2=32'd120;
#400 value1=32'd121;value2=32'd132;
#400 value1=32'd141;value2=32'd157;
#400 value1=32'd159;value2=32'd164;
#400 value1=32'd166;value2=32'd295;
#400 value1=32'd350;value2=32'd395;
#400 value1=32'd441;value2=32'd443;
#400 value1=32'd4;value2=32'd61;
#400 value1=32'd108;value2=32'd110;
#400 value1=32'd122;value2=32'd133;
#400 value1=32'd153;value2=32'd154;
#400 value1=32'd156;value2=32'd157;
#400 value1=32'd160;value2=32'd171;
#400 value1=32'd173;value2=32'd296;
#400 value1=32'd351;value2=32'd396;
#400 value1=32'd448;value2=32'd450;
#400 value1=32'd62;value2=32'd111;
#400 value1=32'd120;value2=32'd123;
#400 value1=32'd134;value2=32'd152;
#400 value1=32'd155;value2=32'd156;
#400 value1=32'd157;value2=32'd161;
#400 value1=32'd177;value2=32'd179;
#400 value1=32'd297;value2=32'd352;
#400 value1=32'd397;value2=32'd456;
#400 value1=32'd4;value2=32'd63;
#400 value1=32'd108;value2=32'd112;
#400 value1=32'd124;value2=32'd135;
#400 value1=32'd152;value2=32'd155;
#400 value1=32'd158;value2=32'd159;
#400 value1=32'd162;value2=32'd182;
#400 value1=32'd184;value2=32'd298;
#400 value1=32'd353;value2=32'd398;
#400 value1=32'd455;value2=32'd461;
#400 value1=32'd64;value2=32'd113;
#400 value1=32'd120;value2=32'd125;
#400 value1=32'd136;value2=32'd153;
#400 value1=32'd154;value2=32'd158;
#400 value1=32'd159;value2=32'd163;
#400 value1=32'd186;value2=32'd188;
#400 value1=32'd299;value2=32'd354;
#400 value1=32'd399;value2=32'd456;
#400 value1=32'd65;value2=32'd114;
#400 value1=32'd126;value2=32'd131;
#400 value1=32'd137;value2=32'd152;
#400 value1=32'd153;value2=32'd157;
#400 value1=32'd158;value2=32'd164;
#400 value1=32'd191;value2=32'd300;
#400 value1=32'd355;value2=32'd400;
#400 value1=32'd457;value2=32'd466;
#400 value1=32'd66;value2=32'd115;
#400 value1=32'd127;value2=32'd138;
#400 value1=32'd141;value2=32'd151;
#400 value1=32'd152;value2=32'd153;
#400 value1=32'd156;value2=32'd159;
#400 value1=32'd165;value2=32'd190;
#400 value1=32'd193;value2=32'd301;
#400 value1=32'd356;value2=32'd401;
#400 value1=32'd458;value2=32'd467;
#400 value1=32'd67;value2=32'd116;
#400 value1=32'd128;value2=32'd131;
#400 value1=32'd139;value2=32'd154;
#400 value1=32'd155;value2=32'd156;
#400 value1=32'd159;value2=32'd166;
#400 value1=32'd191;value2=32'd302;
#400 value1=32'd357;value2=32'd402;
#400 value1=32'd459;value2=32'd468;
#400 value1=32'd68;value2=32'd117;
#400 value1=32'd129;value2=32'd140;
#400 value1=32'd141;value2=32'd151;
#400 value1=32'd154;value2=32'd155;
#400 value1=32'd157;value2=32'd158;
#400 value1=32'd167;value2=32'd192;
#400 value1=32'd195;value2=32'd303;
#400 value1=32'd358;value2=32'd403;
#400 value1=32'd460;value2=32'd469;
#400 value1=32'd5;value2=32'd69;
#400 value1=32'd109;value2=32'd110;
#400 value1=32'd122;value2=32'd143;
#400 value1=32'd152;value2=32'd161;
#400 value1=32'd162;value2=32'd164;
#400 value1=32'd165;value2=32'd172;
#400 value1=32'd174;value2=32'd304;
#400 value1=32'd359;value2=32'd404;
#400 value1=32'd476;value2=32'd478;
#400 value1=32'd70;value2=32'd111;
#400 value1=32'd121;value2=32'd123;
#400 value1=32'd144;value2=32'd153;
#400 value1=32'd160;value2=32'd163;
#400 value1=32'd164;value2=32'd165;
#400 value1=32'd178;value2=32'd180;
#400 value1=32'd305;value2=32'd360;
#400 value1=32'd405;value2=32'd484;
#400 value1=32'd5;value2=32'd71;
#400 value1=32'd109;value2=32'd112;
#400 value1=32'd124;value2=32'd145;
#400 value1=32'd154;value2=32'd160;
#400 value1=32'd163;value2=32'd166;
#400 value1=32'd167;value2=32'd183;
#400 value1=32'd185;value2=32'd306;
#400 value1=32'd361;value2=32'd406;
#400 value1=32'd483;value2=32'd489;
#400 value1=32'd72;value2=32'd113;
#400 value1=32'd121;value2=32'd125;
#400 value1=32'd146;value2=32'd155;
#400 value1=32'd161;value2=32'd162;
#400 value1=32'd166;value2=32'd167;
#400 value1=32'd187;value2=32'd189;
#400 value1=32'd307;value2=32'd362;
#400 value1=32'd407;value2=32'd484;
#400 value1=32'd73;value2=32'd114;
#400 value1=32'd126;value2=32'd132;
#400 value1=32'd147;value2=32'd151;
#400 value1=32'd156;value2=32'd160;
#400 value1=32'd161;value2=32'd165;
#400 value1=32'd166;value2=32'd190;
#400 value1=32'd192;value2=32'd308;
#400 value1=32'd363;value2=32'd408;
#400 value1=32'd485;value2=32'd494;
#400 value1=32'd74;value2=32'd115;
#400 value1=32'd127;value2=32'd142;
#400 value1=32'd148;value2=32'd157;
#400 value1=32'd160;value2=32'd161;
#400 value1=32'd164;value2=32'd167;
#400 value1=32'd194;value2=32'd309;
#400 value1=32'd364;value2=32'd409;
#400 value1=32'd486;value2=32'd495;
#400 value1=32'd75;value2=32'd116;
#400 value1=32'd128;value2=32'd132;
#400 value1=32'd149;value2=32'd151;
#400 value1=32'd158;value2=32'd162;
#400 value1=32'd163;value2=32'd164;
#400 value1=32'd167;value2=32'd193;
#400 value1=32'd195;value2=32'd310;
#400 value1=32'd365;value2=32'd410;
#400 value1=32'd487;value2=32'd496;
#400 value1=32'd76;value2=32'd117;
#400 value1=32'd129;value2=32'd142;
#400 value1=32'd150;value2=32'd159;
#400 value1=32'd162;value2=32'd163;
#400 value1=32'd165;value2=32'd166;
#400 value1=32'd194;value2=32'd311;
#400 value1=32'd366;value2=32'd411;
#400 value1=32'd488;value2=32'd497;
#400 value1=32'd7;value2=32'd77;
#400 value1=32'd111;value2=32'd122;
#400 value1=32'd170;value2=32'd171;
#400 value1=32'd172;value2=32'd175;
#400 value1=32'd177;value2=32'd178;
#400 value1=32'd312;value2=32'd367;
#400 value1=32'd412;value2=32'd505;
#400 value1=32'd6;value2=32'd8;
#400 value1=32'd78;value2=32'd110;
#400 value1=32'd112;value2=32'd170;
#400 value1=32'd173;value2=32'd174;
#400 value1=32'd175;value2=32'd182;
#400 value1=32'd183;value2=32'd313;
#400 value1=32'd368;value2=32'd413;
#400 value1=32'd504;value2=32'd510;
#400 value1=32'd9;value2=32'd79;
#400 value1=32'd113;value2=32'd122;
#400 value1=32'd168;value2=32'd169;
#400 value1=32'd173;value2=32'd174;
#400 value1=32'd176;value2=32'd181;
#400 value1=32'd186;value2=32'd187;
#400 value1=32'd314;value2=32'd369;
#400 value1=32'd414;value2=32'd505;
#400 value1=32'd10;value2=32'd80;
#400 value1=32'd114;value2=32'd133;
#400 value1=32'd152;value2=32'd168;
#400 value1=32'd172;value2=32'd173;
#400 value1=32'd177;value2=32'd182;
#400 value1=32'd190;value2=32'd315;
#400 value1=32'd370;value2=32'd415;
#400 value1=32'd506;value2=32'd515;
#400 value1=32'd11;value2=32'd81;
#400 value1=32'd115;value2=32'd143;
#400 value1=32'd160;value2=32'd168;
#400 value1=32'd171;value2=32'd174;
#400 value1=32'd178;value2=32'd183;
#400 value1=32'd190;value2=32'd316;
#400 value1=32'd371;value2=32'd416;
#400 value1=32'd507;value2=32'd516;
#400 value1=32'd12;value2=32'd82;
#400 value1=32'd116;value2=32'd133;
#400 value1=32'd152;value2=32'd169;
#400 value1=32'd170;value2=32'd171;
#400 value1=32'd174;value2=32'd179;
#400 value1=32'd184;value2=32'd191;
#400 value1=32'd193;value2=32'd317;
#400 value1=32'd372;value2=32'd417;
#400 value1=32'd508;value2=32'd517;
#400 value1=32'd13;value2=32'd83;
#400 value1=32'd117;value2=32'd143;
#400 value1=32'd160;value2=32'd169;
#400 value1=32'd170;value2=32'd172;
#400 value1=32'd173;value2=32'd180;
#400 value1=32'd185;value2=32'd192;
#400 value1=32'd194;value2=32'd318;
#400 value1=32'd373;value2=32'd418;
#400 value1=32'd509;value2=32'd518;
#400 value1=32'd7;value2=32'd84;
#400 value1=32'd111;value2=32'd124;
#400 value1=32'd168;value2=32'd169;
#400 value1=32'd176;value2=32'd179;
#400 value1=32'd180;value2=32'd181;
#400 value1=32'd182;value2=32'd183;
#400 value1=32'd319;value2=32'd374;
#400 value1=32'd419;value2=32'd525;
#400 value1=32'd85;value2=32'd123;
#400 value1=32'd125;value2=32'd170;
#400 value1=32'd175;value2=32'd179;
#400 value1=32'd180;value2=32'd186;
#400 value1=32'd187;value2=32'd320;
#400 value1=32'd375;value2=32'd420;
#400 value1=32'd86;value2=32'd126;
#400 value1=32'd134;value2=32'd153;
#400 value1=32'd168;value2=32'd171;
#400 value1=32'd178;value2=32'd179;
#400 value1=32'd186;value2=32'd190;
#400 value1=32'd321;value2=32'd376;
#400 value1=32'd421;value2=32'd530;
#400 value1=32'd87;value2=32'd127;
#400 value1=32'd144;value2=32'd161;
#400 value1=32'd168;value2=32'd172;
#400 value1=32'd177;value2=32'd180;
#400 value1=32'd187;value2=32'd190;
#400 value1=32'd322;value2=32'd377;
#400 value1=32'd422;value2=32'd531;
#400 value1=32'd88;value2=32'd128;
#400 value1=32'd134;value2=32'd153;
#400 value1=32'd173;value2=32'd175;
#400 value1=32'd176;value2=32'd177;
#400 value1=32'd180;value2=32'd188;
#400 value1=32'd191;value2=32'd193;
#400 value1=32'd323;value2=32'd378;
#400 value1=32'd423;value2=32'd532;
#400 value1=32'd89;value2=32'd129;
#400 value1=32'd144;value2=32'd161;
#400 value1=32'd174;value2=32'd175;
#400 value1=32'd176;value2=32'd178;
#400 value1=32'd179;value2=32'd189;
#400 value1=32'd192;value2=32'd194;
#400 value1=32'd324;value2=32'd379;
#400 value1=32'd424;value2=32'd533;
#400 value1=32'd9;value2=32'd90;
#400 value1=32'd113;value2=32'd124;
#400 value1=32'd170;value2=32'd175;
#400 value1=32'd184;value2=32'd185;
#400 value1=32'd188;value2=32'd189;
#400 value1=32'd325;value2=32'd380;
#400 value1=32'd425;value2=32'd525;
#400 value1=32'd10;value2=32'd91;
#400 value1=32'd114;value2=32'd135;
#400 value1=32'd154;value2=32'd169;
#400 value1=32'd171;value2=32'd175;
#400 value1=32'd183;value2=32'd184;
#400 value1=32'd186;value2=32'd191;
#400 value1=32'd192;value2=32'd326;
#400 value1=32'd381;value2=32'd426;
#400 value1=32'd526;value2=32'd540;
#400 value1=32'd11;value2=32'd92;
#400 value1=32'd115;value2=32'd145;
#400 value1=32'd162;value2=32'd169;
#400 value1=32'd172;value2=32'd175;
#400 value1=32'd182;value2=32'd185;
#400 value1=32'd187;value2=32'd193;
#400 value1=32'd194;value2=32'd327;
#400 value1=32'd382;value2=32'd427;
#400 value1=32'd527;value2=32'd541;
#400 value1=32'd12;value2=32'd93;
#400 value1=32'd116;value2=32'd135;
#400 value1=32'd154;value2=32'd173;
#400 value1=32'd181;value2=32'd182;
#400 value1=32'd185;value2=32'd188;
#400 value1=32'd195;value2=32'd328;
#400 value1=32'd383;value2=32'd428;
#400 value1=32'd528;value2=32'd542;
#400 value1=32'd13;value2=32'd94;
#400 value1=32'd117;value2=32'd145;
#400 value1=32'd162;value2=32'd174;
#400 value1=32'd181;value2=32'd183;
#400 value1=32'd184;value2=32'd189;
#400 value1=32'd195;value2=32'd329;
#400 value1=32'd384;value2=32'd429;
#400 value1=32'd529;value2=32'd543;
#400 value1=32'd95;value2=32'd126;
#400 value1=32'd136;value2=32'd155;
#400 value1=32'd170;value2=32'd176;
#400 value1=32'd177;value2=32'd182;
#400 value1=32'd187;value2=32'd188;
#400 value1=32'd191;value2=32'd192;
#400 value1=32'd330;value2=32'd385;
#400 value1=32'd430;value2=32'd530;
#400 value1=32'd96;value2=32'd127;
#400 value1=32'd146;value2=32'd163;
#400 value1=32'd170;value2=32'd176;
#400 value1=32'd178;value2=32'd183;
#400 value1=32'd186;value2=32'd189;
#400 value1=32'd193;value2=32'd194;
#400 value1=32'd331;value2=32'd386;
#400 value1=32'd431;value2=32'd531;
#400 value1=32'd97;value2=32'd128;
#400 value1=32'd136;value2=32'd155;
#400 value1=32'd179;value2=32'd181;
#400 value1=32'd184;value2=32'd186;
#400 value1=32'd189;value2=32'd195;
#400 value1=32'd332;value2=32'd387;
#400 value1=32'd432;value2=32'd532;
#400 value1=32'd98;value2=32'd129;
#400 value1=32'd146;value2=32'd163;
#400 value1=32'd180;value2=32'd181;
#400 value1=32'd185;value2=32'd187;
#400 value1=32'd188;value2=32'd195;
#400 value1=32'd333;value2=32'd388;
#400 value1=32'd433;value2=32'd533;
#400 value1=32'd99;value2=32'd138;
#400 value1=32'd147;value2=32'd157;
#400 value1=32'd164;value2=32'd171;
#400 value1=32'd172;value2=32'd177;
#400 value1=32'd178;value2=32'd192;
#400 value1=32'd193;value2=32'd334;
#400 value1=32'd389;value2=32'd434;
#400 value1=32'd534;value2=32'd550;
#400 value1=32'd100;value2=32'd137;
#400 value1=32'd139;value2=32'd156;
#400 value1=32'd158;value2=32'd173;
#400 value1=32'd179;value2=32'd182;
#400 value1=32'd186;value2=32'd192;
#400 value1=32'd193;value2=32'd335;
#400 value1=32'd390;value2=32'd435;
#400 value1=32'd535;value2=32'd551;
#400 value1=32'd101;value2=32'd140;
#400 value1=32'd147;value2=32'd159;
#400 value1=32'd164;value2=32'd174;
#400 value1=32'd180;value2=32'd182;
#400 value1=32'd186;value2=32'd190;
#400 value1=32'd191;value2=32'd194;
#400 value1=32'd195;value2=32'd336;
#400 value1=32'd391;value2=32'd436;
#400 value1=32'd536;value2=32'd552;
#400 value1=32'd102;value2=32'd138;
#400 value1=32'd149;value2=32'd157;
#400 value1=32'd166;value2=32'd173;
#400 value1=32'd179;value2=32'd183;
#400 value1=32'd187;value2=32'd190;
#400 value1=32'd191;value2=32'd194;
#400 value1=32'd195;value2=32'd337;
#400 value1=32'd392;value2=32'd437;
#400 value1=32'd537;value2=32'd553;
#400 value1=32'd103;value2=32'd148;
#400 value1=32'd150;value2=32'd165;
#400 value1=32'd167;value2=32'd174;
#400 value1=32'd180;value2=32'd183;
#400 value1=32'd187;value2=32'd192;
#400 value1=32'd193;value2=32'd338;
#400 value1=32'd393;value2=32'd438;
#400 value1=32'd538;value2=32'd554;
#400 value1=32'd104;value2=32'd140;
#400 value1=32'd149;value2=32'd159;
#400 value1=32'd166;value2=32'd184;
#400 value1=32'd185;value2=32'd188;
#400 value1=32'd189;value2=32'd192;
#400 value1=32'd193;value2=32'd339;
#400 value1=32'd394;value2=32'd439;
#400 value1=32'd539;value2=32'd555;
#400 value1=32'd14;value2=32'd27;
#400 value1=32'd105;value2=32'd106;
#400 value1=32'd197;value2=32'd198;
#400 value1=32'd204;value2=32'd206;
#400 value1=32'd209;value2=32'd210;
#400 value1=32'd212;value2=32'd214;
#400 value1=32'd275;value2=32'd276;
#400 value1=32'd277;value2=32'd279;
#400 value1=32'd14;value2=32'd28;
#400 value1=32'd105;value2=32'd107;
#400 value1=32'd196;value2=32'd199;
#400 value1=32'd205;value2=32'd207;
#400 value1=32'd219;value2=32'd220;
#400 value1=32'd222;value2=32'd224;
#400 value1=32'd285;value2=32'd286;
#400 value1=32'd287;value2=32'd289;
#400 value1=32'd29;value2=32'd108;
#400 value1=32'd196;value2=32'd199;
#400 value1=32'd204;value2=32'd206;
#400 value1=32'd229;value2=32'd231;
#400 value1=32'd233;value2=32'd295;
#400 value1=32'd296;value2=32'd298;
#400 value1=32'd30;value2=32'd109;
#400 value1=32'd197;value2=32'd198;
#400 value1=32'd205;value2=32'd207;
#400 value1=32'd229;value2=32'd239;
#400 value1=32'd241;value2=32'd295;
#400 value1=32'd304;value2=32'd306;
#400 value1=32'd14;value2=32'd31;
#400 value1=32'd110;value2=32'd201;
#400 value1=32'd202;value2=32'd204;
#400 value1=32'd205;value2=32'd230;
#400 value1=32'd238;value2=32'd246;
#400 value1=32'd248;value2=32'd296;
#400 value1=32'd304;value2=32'd313;
#400 value1=32'd32;value2=32'd105;
#400 value1=32'd111;value2=32'd200;
#400 value1=32'd203;value2=32'd204;
#400 value1=32'd205;value2=32'd231;
#400 value1=32'd239;value2=32'd254;
#400 value1=32'd297;value2=32'd305;
#400 value1=32'd312;value2=32'd319;
#400 value1=32'd14;value2=32'd33;
#400 value1=32'd112;value2=32'd200;
#400 value1=32'd203;value2=32'd206;
#400 value1=32'd207;value2=32'd232;
#400 value1=32'd240;value2=32'd253;
#400 value1=32'd259;value2=32'd298;
#400 value1=32'd306;value2=32'd313;
#400 value1=32'd34;value2=32'd105;
#400 value1=32'd113;value2=32'd201;
#400 value1=32'd202;value2=32'd206;
#400 value1=32'd207;value2=32'd233;
#400 value1=32'd241;value2=32'd254;
#400 value1=32'd299;value2=32'd307;
#400 value1=32'd314;value2=32'd325;
#400 value1=32'd35;value2=32'd114;
#400 value1=32'd196;value2=32'd198;
#400 value1=32'd200;value2=32'd201;
#400 value1=32'd205;value2=32'd206;
#400 value1=32'd234;value2=32'd242;
#400 value1=32'd255;value2=32'd264;
#400 value1=32'd300;value2=32'd308;
#400 value1=32'd315;value2=32'd326;
#400 value1=32'd36;value2=32'd115;
#400 value1=32'd197;value2=32'd199;
#400 value1=32'd200;value2=32'd201;
#400 value1=32'd204;value2=32'd207;
#400 value1=32'd235;value2=32'd243;
#400 value1=32'd256;value2=32'd265;
#400 value1=32'd301;value2=32'd309;
#400 value1=32'd316;value2=32'd327;
#400 value1=32'd37;value2=32'd116;
#400 value1=32'd196;value2=32'd198;
#400 value1=32'd202;value2=32'd203;
#400 value1=32'd204;value2=32'd207;
#400 value1=32'd236;value2=32'd244;
#400 value1=32'd257;value2=32'd266;
#400 value1=32'd302;value2=32'd310;
#400 value1=32'd317;value2=32'd328;
#400 value1=32'd38;value2=32'd117;
#400 value1=32'd197;value2=32'd199;
#400 value1=32'd202;value2=32'd203;
#400 value1=32'd205;value2=32'd206;
#400 value1=32'd237;value2=32'd245;
#400 value1=32'd258;value2=32'd267;
#400 value1=32'd303;value2=32'd311;
#400 value1=32'd318;value2=32'd329;
#400 value1=32'd15;value2=32'd16;
#400 value1=32'd39;value2=32'd106;
#400 value1=32'd107;value2=32'd210;
#400 value1=32'd216;value2=32'd218;
#400 value1=32'd219;value2=32'd225;
#400 value1=32'd227;value2=32'd274;
#400 value1=32'd340;value2=32'd341;
#400 value1=32'd342;value2=32'd344;
#400 value1=32'd17;value2=32'd40;
#400 value1=32'd108;value2=32'd196;
#400 value1=32'd210;value2=32'd215;
#400 value1=32'd217;value2=32'd219;
#400 value1=32'd234;value2=32'd236;
#400 value1=32'd275;value2=32'd350;
#400 value1=32'd351;value2=32'd353;
#400 value1=32'd18;value2=32'd41;
#400 value1=32'd109;value2=32'd196;
#400 value1=32'd208;value2=32'd209;
#400 value1=32'd216;value2=32'd218;
#400 value1=32'd220;value2=32'd229;
#400 value1=32'd242;value2=32'd244;
#400 value1=32'd276;value2=32'd350;
#400 value1=32'd359;value2=32'd361;
#400 value1=32'd15;value2=32'd19;
#400 value1=32'd42;value2=32'd110;
#400 value1=32'd212;value2=32'd213;
#400 value1=32'd215;value2=32'd216;
#400 value1=32'd221;value2=32'd230;
#400 value1=32'd249;value2=32'd251;
#400 value1=32'd277;value2=32'd351;
#400 value1=32'd359;value2=32'd368;
#400 value1=32'd20;value2=32'd43;
#400 value1=32'd106;value2=32'd111;
#400 value1=32'd196;value2=32'd211;
#400 value1=32'd214;value2=32'd215;
#400 value1=32'd216;value2=32'd222;
#400 value1=32'd231;value2=32'd255;
#400 value1=32'd257;value2=32'd278;
#400 value1=32'd352;value2=32'd360;
#400 value1=32'd367;value2=32'd374;
#400 value1=32'd15;value2=32'd21;
#400 value1=32'd44;value2=32'd112;
#400 value1=32'd211;value2=32'd214;
#400 value1=32'd217;value2=32'd218;
#400 value1=32'd223;value2=32'd232;
#400 value1=32'd260;value2=32'd262;
#400 value1=32'd279;value2=32'd353;
#400 value1=32'd361;value2=32'd368;
#400 value1=32'd22;value2=32'd45;
#400 value1=32'd106;value2=32'd113;
#400 value1=32'd196;value2=32'd212;
#400 value1=32'd213;value2=32'd217;
#400 value1=32'd218;value2=32'd224;
#400 value1=32'd233;value2=32'd264;
#400 value1=32'd266;value2=32'd280;
#400 value1=32'd354;value2=32'd362;
#400 value1=32'd369;value2=32'd380;
#400 value1=32'd23;value2=32'd46;
#400 value1=32'd114;value2=32'd209;
#400 value1=32'd211;value2=32'd212;
#400 value1=32'd216;value2=32'd217;
#400 value1=32'd225;value2=32'd234;
#400 value1=32'd269;value2=32'd281;
#400 value1=32'd355;value2=32'd363;
#400 value1=32'd370;value2=32'd381;
#400 value1=32'd24;value2=32'd47;
#400 value1=32'd115;value2=32'd208;
#400 value1=32'd210;value2=32'd211;
#400 value1=32'd212;value2=32'd215;
#400 value1=32'd218;value2=32'd226;
#400 value1=32'd235;value2=32'd268;
#400 value1=32'd271;value2=32'd282;
#400 value1=32'd356;value2=32'd364;
#400 value1=32'd371;value2=32'd382;
#400 value1=32'd25;value2=32'd48;
#400 value1=32'd116;value2=32'd209;
#400 value1=32'd213;value2=32'd214;
#400 value1=32'd215;value2=32'd218;
#400 value1=32'd227;value2=32'd236;
#400 value1=32'd269;value2=32'd283;
#400 value1=32'd357;value2=32'd365;
#400 value1=32'd372;value2=32'd383;
#400 value1=32'd26;value2=32'd49;
#400 value1=32'd117;value2=32'd208;
#400 value1=32'd210;value2=32'd213;
#400 value1=32'd214;value2=32'd216;
#400 value1=32'd217;value2=32'd228;
#400 value1=32'd237;value2=32'd270;
#400 value1=32'd273;value2=32'd284;
#400 value1=32'd358;value2=32'd366;
#400 value1=32'd373;value2=32'd384;
#400 value1=32'd17;value2=32'd50;
#400 value1=32'd108;value2=32'd197;
#400 value1=32'd208;value2=32'd209;
#400 value1=32'd220;value2=32'd225;
#400 value1=32'd227;value2=32'd229;
#400 value1=32'd235;value2=32'd237;
#400 value1=32'd285;value2=32'd395;
#400 value1=32'd396;value2=32'd398;
#400 value1=32'd18;value2=32'd51;
#400 value1=32'd109;value2=32'd197;
#400 value1=32'd210;value2=32'd219;
#400 value1=32'd226;value2=32'd228;
#400 value1=32'd243;value2=32'd245;
#400 value1=32'd286;value2=32'd395;
#400 value1=32'd404;value2=32'd406;
#400 value1=32'd16;value2=32'd19;
#400 value1=32'd52;value2=32'd110;
#400 value1=32'd211;value2=32'd222;
#400 value1=32'd223;value2=32'd225;
#400 value1=32'd226;value2=32'd238;
#400 value1=32'd250;value2=32'd252;
#400 value1=32'd287;value2=32'd396;
#400 value1=32'd404;value2=32'd413;
#400 value1=32'd20;value2=32'd53;
#400 value1=32'd107;value2=32'd111;
#400 value1=32'd197;value2=32'd212;
#400 value1=32'd221;value2=32'd224;
#400 value1=32'd225;value2=32'd226;
#400 value1=32'd239;value2=32'd256;
#400 value1=32'd258;value2=32'd288;
#400 value1=32'd397;value2=32'd405;
#400 value1=32'd412;value2=32'd419;
#400 value1=32'd16;value2=32'd21;
#400 value1=32'd54;value2=32'd112;
#400 value1=32'd213;value2=32'd221;
#400 value1=32'd224;value2=32'd227;
#400 value1=32'd228;value2=32'd240;
#400 value1=32'd261;value2=32'd263;
#400 value1=32'd289;value2=32'd398;
#400 value1=32'd406;value2=32'd413;
#400 value1=32'd22;value2=32'd55;
#400 value1=32'd107;value2=32'd113;
#400 value1=32'd197;value2=32'd214;
#400 value1=32'd222;value2=32'd223;
#400 value1=32'd227;value2=32'd228;
#400 value1=32'd241;value2=32'd265;
#400 value1=32'd267;value2=32'd290;
#400 value1=32'd399;value2=32'd407;
#400 value1=32'd414;value2=32'd425;
#400 value1=32'd23;value2=32'd56;
#400 value1=32'd114;value2=32'd208;
#400 value1=32'd215;value2=32'd219;
#400 value1=32'd221;value2=32'd222;
#400 value1=32'd226;value2=32'd227;
#400 value1=32'd242;value2=32'd268;
#400 value1=32'd270;value2=32'd291;
#400 value1=32'd400;value2=32'd408;
#400 value1=32'd415;value2=32'd426;
#400 value1=32'd24;value2=32'd57;
#400 value1=32'd115;value2=32'd216;
#400 value1=32'd220;value2=32'd221;
#400 value1=32'd222;value2=32'd225;
#400 value1=32'd228;value2=32'd243;
#400 value1=32'd272;value2=32'd292;
#400 value1=32'd401;value2=32'd409;
#400 value1=32'd416;value2=32'd427;
#400 value1=32'd25;value2=32'd58;
#400 value1=32'd116;value2=32'd208;
#400 value1=32'd217;value2=32'd219;
#400 value1=32'd223;value2=32'd224;
#400 value1=32'd225;value2=32'd228;
#400 value1=32'd244;value2=32'd271;
#400 value1=32'd273;value2=32'd293;
#400 value1=32'd402;value2=32'd410;
#400 value1=32'd417;value2=32'd428;
#400 value1=32'd26;value2=32'd59;
#400 value1=32'd117;value2=32'd218;
#400 value1=32'd220;value2=32'd223;
#400 value1=32'd224;value2=32'd226;
#400 value1=32'd227;value2=32'd245;
#400 value1=32'd272;value2=32'd294;
#400 value1=32'd403;value2=32'd411;
#400 value1=32'd418;value2=32'd429;
#400 value1=32'd60;value2=32'd198;
#400 value1=32'd199;value2=32'd210;
#400 value1=32'd219;value2=32'd235;
#400 value1=32'd237;value2=32'd242;
#400 value1=32'd244;value2=32'd295;
#400 value1=32'd440;value2=32'd442;
#400 value1=32'd17;value2=32'd61;
#400 value1=32'd200;value2=32'd211;
#400 value1=32'd231;value2=32'd232;
#400 value1=32'd234;value2=32'd235;
#400 value1=32'd238;value2=32'd249;
#400 value1=32'd251;value2=32'd296;
#400 value1=32'd440;value2=32'd449;
#400 value1=32'd62;value2=32'd108;
#400 value1=32'd198;value2=32'd201;
#400 value1=32'd212;value2=32'd230;
#400 value1=32'd233;value2=32'd234;
#400 value1=32'd235;value2=32'd239;
#400 value1=32'd255;value2=32'd257;
#400 value1=32'd297;value2=32'd441;
#400 value1=32'd448;value2=32'd455;
#400 value1=32'd17;value2=32'd63;
#400 value1=32'd202;value2=32'd213;
#400 value1=32'd230;value2=32'd233;
#400 value1=32'd236;value2=32'd237;
#400 value1=32'd240;value2=32'd260;
#400 value1=32'd262;value2=32'd298;
#400 value1=32'd442;value2=32'd449;
#400 value1=32'd64;value2=32'd108;
#400 value1=32'd198;value2=32'd203;
#400 value1=32'd214;value2=32'd231;
#400 value1=32'd232;value2=32'd236;
#400 value1=32'd237;value2=32'd241;
#400 value1=32'd264;value2=32'd266;
#400 value1=32'd299;value2=32'd443;
#400 value1=32'd450;value2=32'd461;
#400 value1=32'd65;value2=32'd204;
#400 value1=32'd209;value2=32'd215;
#400 value1=32'd230;value2=32'd231;
#400 value1=32'd235;value2=32'd236;
#400 value1=32'd242;value2=32'd269;
#400 value1=32'd300;value2=32'd444;
#400 value1=32'd451;value2=32'd462;
#400 value1=32'd66;value2=32'd205;
#400 value1=32'd216;value2=32'd219;
#400 value1=32'd229;value2=32'd230;
#400 value1=32'd231;value2=32'd234;
#400 value1=32'd237;value2=32'd243;
#400 value1=32'd268;value2=32'd271;
#400 value1=32'd301;value2=32'd445;
#400 value1=32'd452;value2=32'd463;
#400 value1=32'd67;value2=32'd206;
#400 value1=32'd209;value2=32'd217;
#400 value1=32'd232;value2=32'd233;
#400 value1=32'd234;value2=32'd237;
#400 value1=32'd244;value2=32'd269;
#400 value1=32'd302;value2=32'd446;
#400 value1=32'd453;value2=32'd464;
#400 value1=32'd68;value2=32'd207;
#400 value1=32'd218;value2=32'd219;
#400 value1=32'd229;value2=32'd232;
#400 value1=32'd233;value2=32'd235;
#400 value1=32'd236;value2=32'd245;
#400 value1=32'd270;value2=32'd273;
#400 value1=32'd303;value2=32'd447;
#400 value1=32'd454;value2=32'd465;
#400 value1=32'd18;value2=32'd69;
#400 value1=32'd200;value2=32'd221;
#400 value1=32'd230;value2=32'd239;
#400 value1=32'd240;value2=32'd242;
#400 value1=32'd243;value2=32'd250;
#400 value1=32'd252;value2=32'd304;
#400 value1=32'd440;value2=32'd477;
#400 value1=32'd70;value2=32'd109;
#400 value1=32'd199;value2=32'd201;
#400 value1=32'd222;value2=32'd231;
#400 value1=32'd238;value2=32'd241;
#400 value1=32'd242;value2=32'd243;
#400 value1=32'd256;value2=32'd258;
#400 value1=32'd305;value2=32'd441;
#400 value1=32'd476;value2=32'd483;
#400 value1=32'd18;value2=32'd71;
#400 value1=32'd202;value2=32'd223;
#400 value1=32'd232;value2=32'd238;
#400 value1=32'd241;value2=32'd244;
#400 value1=32'd245;value2=32'd261;
#400 value1=32'd263;value2=32'd306;
#400 value1=32'd442;value2=32'd477;
#400 value1=32'd72;value2=32'd109;
#400 value1=32'd199;value2=32'd203;
#400 value1=32'd224;value2=32'd233;
#400 value1=32'd239;value2=32'd240;
#400 value1=32'd244;value2=32'd245;
#400 value1=32'd265;value2=32'd267;
#400 value1=32'd307;value2=32'd443;
#400 value1=32'd478;value2=32'd489;
#400 value1=32'd73;value2=32'd204;
#400 value1=32'd210;value2=32'd225;
#400 value1=32'd229;value2=32'd234;
#400 value1=32'd238;value2=32'd239;
#400 value1=32'd243;value2=32'd244;
#400 value1=32'd268;value2=32'd270;
#400 value1=32'd308;value2=32'd444;
#400 value1=32'd479;value2=32'd490;
#400 value1=32'd74;value2=32'd205;
#400 value1=32'd220;value2=32'd226;
#400 value1=32'd235;value2=32'd238;
#400 value1=32'd239;value2=32'd242;
#400 value1=32'd245;value2=32'd272;
#400 value1=32'd309;value2=32'd445;
#400 value1=32'd480;value2=32'd491;
#400 value1=32'd75;value2=32'd206;
#400 value1=32'd210;value2=32'd227;
#400 value1=32'd229;value2=32'd236;
#400 value1=32'd240;value2=32'd241;
#400 value1=32'd242;value2=32'd245;
#400 value1=32'd271;value2=32'd273;
#400 value1=32'd310;value2=32'd446;
#400 value1=32'd481;value2=32'd492;
#400 value1=32'd76;value2=32'd207;
#400 value1=32'd220;value2=32'd228;
#400 value1=32'd237;value2=32'd240;
#400 value1=32'd241;value2=32'd243;
#400 value1=32'd244;value2=32'd272;
#400 value1=32'd311;value2=32'd447;
#400 value1=32'd482;value2=32'd493;
#400 value1=32'd20;value2=32'd77;
#400 value1=32'd110;value2=32'd200;
#400 value1=32'd248;value2=32'd249;
#400 value1=32'd250;value2=32'd253;
#400 value1=32'd255;value2=32'd256;
#400 value1=32'd312;value2=32'd448;
#400 value1=32'd476;value2=32'd504;
#400 value1=32'd19;value2=32'd21;
#400 value1=32'd78;value2=32'd248;
#400 value1=32'd251;value2=32'd252;
#400 value1=32'd253;value2=32'd260;
#400 value1=32'd261;value2=32'd313;
#400 value1=32'd449;value2=32'd477;
#400 value1=32'd22;value2=32'd79;
#400 value1=32'd110;value2=32'd200;
#400 value1=32'd246;value2=32'd247;
#400 value1=32'd251;value2=32'd252;
#400 value1=32'd254;value2=32'd259;
#400 value1=32'd264;value2=32'd265;
#400 value1=32'd314;value2=32'd450;
#400 value1=32'd478;value2=32'd510;
#400 value1=32'd23;value2=32'd80;
#400 value1=32'd211;value2=32'd230;
#400 value1=32'd246;value2=32'd250;
#400 value1=32'd251;value2=32'd255;
#400 value1=32'd260;value2=32'd268;
#400 value1=32'd315;value2=32'd451;
#400 value1=32'd479;value2=32'd511;
#400 value1=32'd24;value2=32'd81;
#400 value1=32'd221;value2=32'd238;
#400 value1=32'd246;value2=32'd249;
#400 value1=32'd252;value2=32'd256;
#400 value1=32'd261;value2=32'd268;
#400 value1=32'd316;value2=32'd452;
#400 value1=32'd480;value2=32'd512;
#400 value1=32'd25;value2=32'd82;
#400 value1=32'd211;value2=32'd230;
#400 value1=32'd247;value2=32'd248;
#400 value1=32'd249;value2=32'd252;
#400 value1=32'd257;value2=32'd262;
#400 value1=32'd269;value2=32'd271;
#400 value1=32'd317;value2=32'd453;
#400 value1=32'd481;value2=32'd513;
#400 value1=32'd26;value2=32'd83;
#400 value1=32'd221;value2=32'd238;
#400 value1=32'd247;value2=32'd248;
#400 value1=32'd250;value2=32'd251;
#400 value1=32'd258;value2=32'd263;
#400 value1=32'd270;value2=32'd272;
#400 value1=32'd318;value2=32'd454;
#400 value1=32'd482;value2=32'd514;
#400 value1=32'd20;value2=32'd84;
#400 value1=32'd112;value2=32'd202;
#400 value1=32'd246;value2=32'd247;
#400 value1=32'd254;value2=32'd257;
#400 value1=32'd258;value2=32'd259;
#400 value1=32'd260;value2=32'd261;
#400 value1=32'd319;value2=32'd455;
#400 value1=32'd483;value2=32'd504;
#400 value1=32'd85;value2=32'd111;
#400 value1=32'd113;value2=32'd201;
#400 value1=32'd203;value2=32'd248;
#400 value1=32'd253;value2=32'd257;
#400 value1=32'd258;value2=32'd264;
#400 value1=32'd265;value2=32'd320;
#400 value1=32'd456;value2=32'd484;
#400 value1=32'd505;value2=32'd525;
#400 value1=32'd86;value2=32'd114;
#400 value1=32'd204;value2=32'd212;
#400 value1=32'd231;value2=32'd246;
#400 value1=32'd249;value2=32'd256;
#400 value1=32'd257;value2=32'd264;
#400 value1=32'd268;value2=32'd321;
#400 value1=32'd457;value2=32'd485;
#400 value1=32'd506;value2=32'd526;
#400 value1=32'd87;value2=32'd115;
#400 value1=32'd205;value2=32'd222;
#400 value1=32'd239;value2=32'd246;
#400 value1=32'd250;value2=32'd255;
#400 value1=32'd258;value2=32'd265;
#400 value1=32'd268;value2=32'd322;
#400 value1=32'd458;value2=32'd486;
#400 value1=32'd507;value2=32'd527;
#400 value1=32'd88;value2=32'd116;
#400 value1=32'd206;value2=32'd212;
#400 value1=32'd231;value2=32'd251;
#400 value1=32'd253;value2=32'd254;
#400 value1=32'd255;value2=32'd258;
#400 value1=32'd266;value2=32'd269;
#400 value1=32'd271;value2=32'd323;
#400 value1=32'd459;value2=32'd487;
#400 value1=32'd508;value2=32'd528;
#400 value1=32'd89;value2=32'd117;
#400 value1=32'd207;value2=32'd222;
#400 value1=32'd239;value2=32'd252;
#400 value1=32'd253;value2=32'd254;
#400 value1=32'd256;value2=32'd257;
#400 value1=32'd267;value2=32'd270;
#400 value1=32'd272;value2=32'd324;
#400 value1=32'd460;value2=32'd488;
#400 value1=32'd509;value2=32'd529;
#400 value1=32'd22;value2=32'd90;
#400 value1=32'd112;value2=32'd202;
#400 value1=32'd248;value2=32'd253;
#400 value1=32'd262;value2=32'd263;
#400 value1=32'd266;value2=32'd267;
#400 value1=32'd325;value2=32'd461;
#400 value1=32'd489;value2=32'd510;
#400 value1=32'd23;value2=32'd91;
#400 value1=32'd213;value2=32'd232;
#400 value1=32'd247;value2=32'd249;
#400 value1=32'd253;value2=32'd261;
#400 value1=32'd262;value2=32'd264;
#400 value1=32'd269;value2=32'd270;
#400 value1=32'd326;value2=32'd462;
#400 value1=32'd490;value2=32'd511;
#400 value1=32'd24;value2=32'd92;
#400 value1=32'd223;value2=32'd240;
#400 value1=32'd247;value2=32'd250;
#400 value1=32'd253;value2=32'd260;
#400 value1=32'd263;value2=32'd265;
#400 value1=32'd271;value2=32'd272;
#400 value1=32'd327;value2=32'd463;
#400 value1=32'd491;value2=32'd512;
#400 value1=32'd25;value2=32'd93;
#400 value1=32'd213;value2=32'd232;
#400 value1=32'd251;value2=32'd259;
#400 value1=32'd260;value2=32'd263;
#400 value1=32'd266;value2=32'd273;
#400 value1=32'd328;value2=32'd464;
#400 value1=32'd492;value2=32'd513;
#400 value1=32'd26;value2=32'd94;
#400 value1=32'd223;value2=32'd240;
#400 value1=32'd252;value2=32'd259;
#400 value1=32'd261;value2=32'd262;
#400 value1=32'd267;value2=32'd273;
#400 value1=32'd329;value2=32'd465;
#400 value1=32'd493;value2=32'd514;
#400 value1=32'd95;value2=32'd114;
#400 value1=32'd204;value2=32'd214;
#400 value1=32'd233;value2=32'd248;
#400 value1=32'd254;value2=32'd255;
#400 value1=32'd260;value2=32'd265;
#400 value1=32'd266;value2=32'd269;
#400 value1=32'd270;value2=32'd330;
#400 value1=32'd466;value2=32'd494;
#400 value1=32'd515;value2=32'd540;
#400 value1=32'd96;value2=32'd115;
#400 value1=32'd205;value2=32'd224;
#400 value1=32'd241;value2=32'd248;
#400 value1=32'd254;value2=32'd256;
#400 value1=32'd261;value2=32'd264;
#400 value1=32'd267;value2=32'd271;
#400 value1=32'd272;value2=32'd331;
#400 value1=32'd467;value2=32'd495;
#400 value1=32'd516;value2=32'd541;
#400 value1=32'd97;value2=32'd116;
#400 value1=32'd206;value2=32'd214;
#400 value1=32'd233;value2=32'd257;
#400 value1=32'd259;value2=32'd262;
#400 value1=32'd264;value2=32'd267;
#400 value1=32'd273;value2=32'd332;
#400 value1=32'd468;value2=32'd496;
#400 value1=32'd517;value2=32'd542;
#400 value1=32'd98;value2=32'd117;
#400 value1=32'd207;value2=32'd224;
#400 value1=32'd241;value2=32'd258;
#400 value1=32'd259;value2=32'd263;
#400 value1=32'd265;value2=32'd266;
#400 value1=32'd273;value2=32'd333;
#400 value1=32'd469;value2=32'd497;
#400 value1=32'd518;value2=32'd543;
#400 value1=32'd99;value2=32'd216;
#400 value1=32'd225;value2=32'd235;
#400 value1=32'd242;value2=32'd249;
#400 value1=32'd250;value2=32'd255;
#400 value1=32'd256;value2=32'd270;
#400 value1=32'd271;value2=32'd334;
#400 value1=32'd470;value2=32'd498;
#400 value1=32'd519;value2=32'd544;
#400 value1=32'd100;value2=32'd215;
#400 value1=32'd217;value2=32'd234;
#400 value1=32'd236;value2=32'd251;
#400 value1=32'd257;value2=32'd260;
#400 value1=32'd264;value2=32'd270;
#400 value1=32'd271;value2=32'd335;
#400 value1=32'd471;value2=32'd499;
#400 value1=32'd520;value2=32'd545;
#400 value1=32'd101;value2=32'd218;
#400 value1=32'd225;value2=32'd237;
#400 value1=32'd242;value2=32'd252;
#400 value1=32'd258;value2=32'd260;
#400 value1=32'd264;value2=32'd268;
#400 value1=32'd269;value2=32'd272;
#400 value1=32'd273;value2=32'd336;
#400 value1=32'd472;value2=32'd500;
#400 value1=32'd521;value2=32'd546;
#400 value1=32'd102;value2=32'd216;
#400 value1=32'd227;value2=32'd235;
#400 value1=32'd244;value2=32'd251;
#400 value1=32'd257;value2=32'd261;
#400 value1=32'd265;value2=32'd268;
#400 value1=32'd269;value2=32'd272;
#400 value1=32'd273;value2=32'd337;
#400 value1=32'd473;value2=32'd501;
#400 value1=32'd522;value2=32'd547;
#400 value1=32'd103;value2=32'd226;
#400 value1=32'd228;value2=32'd243;
#400 value1=32'd245;value2=32'd252;
#400 value1=32'd258;value2=32'd261;
#400 value1=32'd265;value2=32'd270;
#400 value1=32'd271;value2=32'd338;
#400 value1=32'd474;value2=32'd502;
#400 value1=32'd523;value2=32'd548;
#400 value1=32'd104;value2=32'd218;
#400 value1=32'd227;value2=32'd237;
#400 value1=32'd244;value2=32'd262;
#400 value1=32'd263;value2=32'd266;
#400 value1=32'd267;value2=32'd270;
#400 value1=32'd271;value2=32'd339;
#400 value1=32'd475;value2=32'd503;
#400 value1=32'd524;value2=32'd549;
#400 value1=32'd27;value2=32'd28;
#400 value1=32'd118;value2=32'd119;
#400 value1=32'd130;value2=32'd208;
#400 value1=32'd276;value2=32'd282;
#400 value1=32'd284;value2=32'd285;
#400 value1=32'd291;value2=32'd293;
#400 value1=32'd340;value2=32'd341;
#400 value1=32'd343;value2=32'd345;
#400 value1=32'd29;value2=32'd120;
#400 value1=32'd131;value2=32'd196;
#400 value1=32'd209;value2=32'd276;
#400 value1=32'd281;value2=32'd283;
#400 value1=32'd285;value2=32'd300;
#400 value1=32'd302;value2=32'd350;
#400 value1=32'd352;value2=32'd354;
#400 value1=32'd30;value2=32'd121;
#400 value1=32'd132;value2=32'd196;
#400 value1=32'd210;value2=32'd274;
#400 value1=32'd275;value2=32'd282;
#400 value1=32'd284;value2=32'd286;
#400 value1=32'd295;value2=32'd308;
#400 value1=32'd310;value2=32'd350;
#400 value1=32'd360;value2=32'd362;
#400 value1=32'd27;value2=32'd31;
#400 value1=32'd122;value2=32'd133;
#400 value1=32'd196;value2=32'd211;
#400 value1=32'd278;value2=32'd279;
#400 value1=32'd281;value2=32'd282;
#400 value1=32'd287;value2=32'd296;
#400 value1=32'd315;value2=32'd317;
#400 value1=32'd351;value2=32'd359;
#400 value1=32'd367;value2=32'd369;
#400 value1=32'd32;value2=32'd118;
#400 value1=32'd123;value2=32'd134;
#400 value1=32'd212;value2=32'd277;
#400 value1=32'd280;value2=32'd281;
#400 value1=32'd282;value2=32'd288;
#400 value1=32'd297;value2=32'd321;
#400 value1=32'd323;value2=32'd352;
#400 value1=32'd360;value2=32'd375;
#400 value1=32'd27;value2=32'd33;
#400 value1=32'd124;value2=32'd135;
#400 value1=32'd196;value2=32'd213;
#400 value1=32'd277;value2=32'd280;
#400 value1=32'd283;value2=32'd284;
#400 value1=32'd289;value2=32'd298;
#400 value1=32'd326;value2=32'd328;
#400 value1=32'd353;value2=32'd361;
#400 value1=32'd374;value2=32'd380;
#400 value1=32'd34;value2=32'd118;
#400 value1=32'd125;value2=32'd136;
#400 value1=32'd214;value2=32'd278;
#400 value1=32'd279;value2=32'd283;
#400 value1=32'd284;value2=32'd290;
#400 value1=32'd299;value2=32'd330;
#400 value1=32'd332;value2=32'd354;
#400 value1=32'd362;value2=32'd375;
#400 value1=32'd35;value2=32'd126;
#400 value1=32'd137;value2=32'd215;
#400 value1=32'd275;value2=32'd277;
#400 value1=32'd278;value2=32'd282;
#400 value1=32'd283;value2=32'd291;
#400 value1=32'd300;value2=32'd335;
#400 value1=32'd355;value2=32'd363;
#400 value1=32'd376;value2=32'd385;
#400 value1=32'd36;value2=32'd127;
#400 value1=32'd138;value2=32'd216;
#400 value1=32'd274;value2=32'd276;
#400 value1=32'd277;value2=32'd278;
#400 value1=32'd281;value2=32'd284;
#400 value1=32'd292;value2=32'd301;
#400 value1=32'd334;value2=32'd337;
#400 value1=32'd356;value2=32'd364;
#400 value1=32'd377;value2=32'd386;
#400 value1=32'd37;value2=32'd128;
#400 value1=32'd139;value2=32'd217;
#400 value1=32'd275;value2=32'd279;
#400 value1=32'd280;value2=32'd281;
#400 value1=32'd284;value2=32'd293;
#400 value1=32'd302;value2=32'd335;
#400 value1=32'd357;value2=32'd365;
#400 value1=32'd378;value2=32'd387;
#400 value1=32'd38;value2=32'd129;
#400 value1=32'd140;value2=32'd218;
#400 value1=32'd274;value2=32'd276;
#400 value1=32'd279;value2=32'd280;
#400 value1=32'd282;value2=32'd283;
#400 value1=32'd294;value2=32'd303;
#400 value1=32'd336;value2=32'd339;
#400 value1=32'd358;value2=32'd366;
#400 value1=32'd379;value2=32'd388;
#400 value1=32'd29;value2=32'd120;
#400 value1=32'd141;value2=32'd197;
#400 value1=32'd219;value2=32'd274;
#400 value1=32'd275;value2=32'd286;
#400 value1=32'd291;value2=32'd293;
#400 value1=32'd295;value2=32'd301;
#400 value1=32'd303;value2=32'd395;
#400 value1=32'd397;value2=32'd399;
#400 value1=32'd30;value2=32'd121;
#400 value1=32'd142;value2=32'd197;
#400 value1=32'd220;value2=32'd276;
#400 value1=32'd285;value2=32'd292;
#400 value1=32'd294;value2=32'd309;
#400 value1=32'd311;value2=32'd395;
#400 value1=32'd405;value2=32'd407;
#400 value1=32'd28;value2=32'd31;
#400 value1=32'd122;value2=32'd143;
#400 value1=32'd197;value2=32'd221;
#400 value1=32'd277;value2=32'd288;
#400 value1=32'd289;value2=32'd291;
#400 value1=32'd292;value2=32'd304;
#400 value1=32'd316;value2=32'd318;
#400 value1=32'd396;value2=32'd404;
#400 value1=32'd412;value2=32'd414;
#400 value1=32'd32;value2=32'd119;
#400 value1=32'd123;value2=32'd144;
#400 value1=32'd222;value2=32'd278;
#400 value1=32'd287;value2=32'd290;
#400 value1=32'd291;value2=32'd292;
#400 value1=32'd305;value2=32'd322;
#400 value1=32'd324;value2=32'd397;
#400 value1=32'd405;value2=32'd420;
#400 value1=32'd28;value2=32'd33;
#400 value1=32'd124;value2=32'd145;
#400 value1=32'd197;value2=32'd223;
#400 value1=32'd279;value2=32'd287;
#400 value1=32'd290;value2=32'd293;
#400 value1=32'd294;value2=32'd306;
#400 value1=32'd327;value2=32'd329;
#400 value1=32'd398;value2=32'd406;
#400 value1=32'd419;value2=32'd425;
#400 value1=32'd34;value2=32'd119;
#400 value1=32'd125;value2=32'd146;
#400 value1=32'd224;value2=32'd280;
#400 value1=32'd288;value2=32'd289;
#400 value1=32'd293;value2=32'd294;
#400 value1=32'd307;value2=32'd331;
#400 value1=32'd333;value2=32'd399;
#400 value1=32'd407;value2=32'd420;
#400 value1=32'd35;value2=32'd126;
#400 value1=32'd147;value2=32'd225;
#400 value1=32'd274;value2=32'd281;
#400 value1=32'd285;value2=32'd287;
#400 value1=32'd288;value2=32'd292;
#400 value1=32'd293;value2=32'd308;
#400 value1=32'd334;value2=32'd336;
#400 value1=32'd400;value2=32'd408;
#400 value1=32'd421;value2=32'd430;
#400 value1=32'd36;value2=32'd127;
#400 value1=32'd148;value2=32'd226;
#400 value1=32'd282;value2=32'd286;
#400 value1=32'd287;value2=32'd288;
#400 value1=32'd291;value2=32'd294;
#400 value1=32'd309;value2=32'd338;
#400 value1=32'd401;value2=32'd409;
#400 value1=32'd422;value2=32'd431;
#400 value1=32'd37;value2=32'd128;
#400 value1=32'd149;value2=32'd227;
#400 value1=32'd274;value2=32'd283;
#400 value1=32'd285;value2=32'd289;
#400 value1=32'd290;value2=32'd291;
#400 value1=32'd294;value2=32'd310;
#400 value1=32'd337;value2=32'd339;
#400 value1=32'd402;value2=32'd410;
#400 value1=32'd423;value2=32'd432;
#400 value1=32'd38;value2=32'd129;
#400 value1=32'd150;value2=32'd228;
#400 value1=32'd284;value2=32'd286;
#400 value1=32'd289;value2=32'd290;
#400 value1=32'd292;value2=32'd293;
#400 value1=32'd311;value2=32'd338;
#400 value1=32'd403;value2=32'd411;
#400 value1=32'd424;value2=32'd433;
#400 value1=32'd151;value2=32'd198;
#400 value1=32'd199;value2=32'd229;
#400 value1=32'd276;value2=32'd285;
#400 value1=32'd301;value2=32'd303;
#400 value1=32'd308;value2=32'd310;
#400 value1=32'd441;value2=32'd443;
#400 value1=32'd29;value2=32'd152;
#400 value1=32'd198;value2=32'd200;
#400 value1=32'd230;value2=32'd277;
#400 value1=32'd297;value2=32'd298;
#400 value1=32'd300;value2=32'd301;
#400 value1=32'd304;value2=32'd315;
#400 value1=32'd317;value2=32'd440;
#400 value1=32'd448;value2=32'd450;
#400 value1=32'd120;value2=32'd153;
#400 value1=32'd201;value2=32'd231;
#400 value1=32'd278;value2=32'd296;
#400 value1=32'd299;value2=32'd300;
#400 value1=32'd301;value2=32'd305;
#400 value1=32'd321;value2=32'd323;
#400 value1=32'd441;value2=32'd456;
#400 value1=32'd29;value2=32'd154;
#400 value1=32'd198;value2=32'd202;
#400 value1=32'd232;value2=32'd279;
#400 value1=32'd296;value2=32'd299;
#400 value1=32'd302;value2=32'd303;
#400 value1=32'd306;value2=32'd326;
#400 value1=32'd328;value2=32'd442;
#400 value1=32'd455;value2=32'd461;
#400 value1=32'd120;value2=32'd155;
#400 value1=32'd203;value2=32'd233;
#400 value1=32'd280;value2=32'd297;
#400 value1=32'd298;value2=32'd302;
#400 value1=32'd303;value2=32'd307;
#400 value1=32'd330;value2=32'd332;
#400 value1=32'd443;value2=32'd456;
#400 value1=32'd156;value2=32'd204;
#400 value1=32'd234;value2=32'd275;
#400 value1=32'd281;value2=32'd296;
#400 value1=32'd297;value2=32'd301;
#400 value1=32'd302;value2=32'd308;
#400 value1=32'd335;value2=32'd444;
#400 value1=32'd457;value2=32'd466;
#400 value1=32'd157;value2=32'd205;
#400 value1=32'd235;value2=32'd282;
#400 value1=32'd285;value2=32'd295;
#400 value1=32'd296;value2=32'd297;
#400 value1=32'd300;value2=32'd303;
#400 value1=32'd309;value2=32'd334;
#400 value1=32'd337;value2=32'd445;
#400 value1=32'd458;value2=32'd467;
#400 value1=32'd158;value2=32'd206;
#400 value1=32'd236;value2=32'd275;
#400 value1=32'd283;value2=32'd298;
#400 value1=32'd299;value2=32'd300;
#400 value1=32'd303;value2=32'd310;
#400 value1=32'd335;value2=32'd446;
#400 value1=32'd459;value2=32'd468;
#400 value1=32'd159;value2=32'd207;
#400 value1=32'd237;value2=32'd284;
#400 value1=32'd285;value2=32'd295;
#400 value1=32'd298;value2=32'd299;
#400 value1=32'd301;value2=32'd302;
#400 value1=32'd311;value2=32'd336;
#400 value1=32'd339;value2=32'd447;
#400 value1=32'd460;value2=32'd469;
#400 value1=32'd30;value2=32'd160;
#400 value1=32'd199;value2=32'd200;
#400 value1=32'd238;value2=32'd287;
#400 value1=32'd296;value2=32'd305;
#400 value1=32'd306;value2=32'd308;
#400 value1=32'd309;value2=32'd316;
#400 value1=32'd318;value2=32'd440;
#400 value1=32'd476;value2=32'd478;
#400 value1=32'd121;value2=32'd161;
#400 value1=32'd201;value2=32'd239;
#400 value1=32'd288;value2=32'd297;
#400 value1=32'd304;value2=32'd307;
#400 value1=32'd308;value2=32'd309;
#400 value1=32'd322;value2=32'd324;
#400 value1=32'd441;value2=32'd484;
#400 value1=32'd30;value2=32'd162;
#400 value1=32'd199;value2=32'd202;
#400 value1=32'd240;value2=32'd289;
#400 value1=32'd298;value2=32'd304;
#400 value1=32'd307;value2=32'd310;
#400 value1=32'd311;value2=32'd327;
#400 value1=32'd329;value2=32'd442;
#400 value1=32'd483;value2=32'd489;
#400 value1=32'd121;value2=32'd163;
#400 value1=32'd203;value2=32'd241;
#400 value1=32'd290;value2=32'd299;
#400 value1=32'd305;value2=32'd306;
#400 value1=32'd310;value2=32'd311;
#400 value1=32'd331;value2=32'd333;
#400 value1=32'd443;value2=32'd484;
#400 value1=32'd164;value2=32'd204;
#400 value1=32'd242;value2=32'd276;
#400 value1=32'd291;value2=32'd295;
#400 value1=32'd300;value2=32'd304;
#400 value1=32'd305;value2=32'd309;
#400 value1=32'd310;value2=32'd334;
#400 value1=32'd336;value2=32'd444;
#400 value1=32'd485;value2=32'd494;
#400 value1=32'd165;value2=32'd205;
#400 value1=32'd243;value2=32'd286;
#400 value1=32'd292;value2=32'd301;
#400 value1=32'd304;value2=32'd305;
#400 value1=32'd308;value2=32'd311;
#400 value1=32'd338;value2=32'd445;
#400 value1=32'd486;value2=32'd495;
#400 value1=32'd166;value2=32'd206;
#400 value1=32'd244;value2=32'd276;
#400 value1=32'd293;value2=32'd295;
#400 value1=32'd302;value2=32'd306;
#400 value1=32'd307;value2=32'd308;
#400 value1=32'd311;value2=32'd337;
#400 value1=32'd339;value2=32'd446;
#400 value1=32'd487;value2=32'd496;
#400 value1=32'd167;value2=32'd207;
#400 value1=32'd245;value2=32'd286;
#400 value1=32'd294;value2=32'd303;
#400 value1=32'd306;value2=32'd307;
#400 value1=32'd309;value2=32'd310;
#400 value1=32'd338;value2=32'd447;
#400 value1=32'd488;value2=32'd497;
#400 value1=32'd32;value2=32'd122;
#400 value1=32'd168;value2=32'd201;
#400 value1=32'd246;value2=32'd314;
#400 value1=32'd315;value2=32'd316;
#400 value1=32'd319;value2=32'd321;
#400 value1=32'd322;value2=32'd448;
#400 value1=32'd476;value2=32'd505;
#400 value1=32'd31;value2=32'd33;
#400 value1=32'd169;value2=32'd200;
#400 value1=32'd202;value2=32'd247;
#400 value1=32'd314;value2=32'd317;
#400 value1=32'd318;value2=32'd319;
#400 value1=32'd326;value2=32'd327;
#400 value1=32'd449;value2=32'd477;
#400 value1=32'd504;value2=32'd510;
#400 value1=32'd34;value2=32'd122;
#400 value1=32'd170;value2=32'd203;
#400 value1=32'd248;value2=32'd312;
#400 value1=32'd313;value2=32'd317;
#400 value1=32'd318;value2=32'd320;
#400 value1=32'd325;value2=32'd330;
#400 value1=32'd331;value2=32'd450;
#400 value1=32'd478;value2=32'd505;
#400 value1=32'd35;value2=32'd171;
#400 value1=32'd204;value2=32'd249;
#400 value1=32'd277;value2=32'd296;
#400 value1=32'd312;value2=32'd316;
#400 value1=32'd317;value2=32'd321;
#400 value1=32'd326;value2=32'd334;
#400 value1=32'd451;value2=32'd479;
#400 value1=32'd506;value2=32'd515;
#400 value1=32'd36;value2=32'd172;
#400 value1=32'd205;value2=32'd250;
#400 value1=32'd287;value2=32'd304;
#400 value1=32'd312;value2=32'd315;
#400 value1=32'd318;value2=32'd322;
#400 value1=32'd327;value2=32'd334;
#400 value1=32'd452;value2=32'd480;
#400 value1=32'd507;value2=32'd516;
#400 value1=32'd37;value2=32'd173;
#400 value1=32'd206;value2=32'd251;
#400 value1=32'd277;value2=32'd296;
#400 value1=32'd313;value2=32'd314;
#400 value1=32'd315;value2=32'd318;
#400 value1=32'd323;value2=32'd328;
#400 value1=32'd335;value2=32'd337;
#400 value1=32'd453;value2=32'd481;
#400 value1=32'd508;value2=32'd517;
#400 value1=32'd38;value2=32'd174;
#400 value1=32'd207;value2=32'd252;
#400 value1=32'd287;value2=32'd304;
#400 value1=32'd313;value2=32'd314;
#400 value1=32'd316;value2=32'd317;
#400 value1=32'd324;value2=32'd329;
#400 value1=32'd336;value2=32'd338;
#400 value1=32'd454;value2=32'd482;
#400 value1=32'd509;value2=32'd518;
#400 value1=32'd32;value2=32'd124;
#400 value1=32'd175;value2=32'd201;
#400 value1=32'd253;value2=32'd312;
#400 value1=32'd313;value2=32'd320;
#400 value1=32'd323;value2=32'd324;
#400 value1=32'd325;value2=32'd326;
#400 value1=32'd327;value2=32'd455;
#400 value1=32'd483;value2=32'd525;
#400 value1=32'd123;value2=32'd125;
#400 value1=32'd176;value2=32'd254;
#400 value1=32'd314;value2=32'd319;
#400 value1=32'd323;value2=32'd324;
#400 value1=32'd330;value2=32'd331;
#400 value1=32'd456;value2=32'd484;
#400 value1=32'd126;value2=32'd177;
#400 value1=32'd255;value2=32'd278;
#400 value1=32'd297;value2=32'd312;
#400 value1=32'd315;value2=32'd322;
#400 value1=32'd323;value2=32'd330;
#400 value1=32'd334;value2=32'd457;
#400 value1=32'd485;value2=32'd530;
#400 value1=32'd127;value2=32'd178;
#400 value1=32'd256;value2=32'd288;
#400 value1=32'd305;value2=32'd312;
#400 value1=32'd316;value2=32'd321;
#400 value1=32'd324;value2=32'd331;
#400 value1=32'd334;value2=32'd458;
#400 value1=32'd486;value2=32'd531;
#400 value1=32'd128;value2=32'd179;
#400 value1=32'd257;value2=32'd278;
#400 value1=32'd297;value2=32'd317;
#400 value1=32'd319;value2=32'd320;
#400 value1=32'd321;value2=32'd324;
#400 value1=32'd332;value2=32'd335;
#400 value1=32'd337;value2=32'd459;
#400 value1=32'd487;value2=32'd532;
#400 value1=32'd129;value2=32'd180;
#400 value1=32'd258;value2=32'd288;
#400 value1=32'd305;value2=32'd318;
#400 value1=32'd319;value2=32'd320;
#400 value1=32'd322;value2=32'd323;
#400 value1=32'd333;value2=32'd336;
#400 value1=32'd338;value2=32'd460;
#400 value1=32'd488;value2=32'd533;
#400 value1=32'd34;value2=32'd124;
#400 value1=32'd181;value2=32'd203;
#400 value1=32'd259;value2=32'd314;
#400 value1=32'd319;value2=32'd328;
#400 value1=32'd329;value2=32'd332;
#400 value1=32'd333;value2=32'd461;
#400 value1=32'd489;value2=32'd525;
#400 value1=32'd35;value2=32'd182;
#400 value1=32'd204;value2=32'd260;
#400 value1=32'd279;value2=32'd298;
#400 value1=32'd313;value2=32'd315;
#400 value1=32'd319;value2=32'd327;
#400 value1=32'd328;value2=32'd330;
#400 value1=32'd335;value2=32'd336;
#400 value1=32'd462;value2=32'd490;
#400 value1=32'd526;value2=32'd540;
#400 value1=32'd36;value2=32'd183;
#400 value1=32'd205;value2=32'd261;
#400 value1=32'd289;value2=32'd306;
#400 value1=32'd313;value2=32'd316;
#400 value1=32'd319;value2=32'd326;
#400 value1=32'd329;value2=32'd331;
#400 value1=32'd337;value2=32'd338;
#400 value1=32'd463;value2=32'd491;
#400 value1=32'd527;value2=32'd541;
#400 value1=32'd37;value2=32'd184;
#400 value1=32'd206;value2=32'd262;
#400 value1=32'd279;value2=32'd298;
#400 value1=32'd317;value2=32'd325;
#400 value1=32'd326;value2=32'd329;
#400 value1=32'd332;value2=32'd339;
#400 value1=32'd464;value2=32'd492;
#400 value1=32'd528;value2=32'd542;
#400 value1=32'd38;value2=32'd185;
#400 value1=32'd207;value2=32'd263;
#400 value1=32'd289;value2=32'd306;
#400 value1=32'd318;value2=32'd325;
#400 value1=32'd327;value2=32'd328;
#400 value1=32'd333;value2=32'd339;
#400 value1=32'd465;value2=32'd493;
#400 value1=32'd529;value2=32'd543;
#400 value1=32'd126;value2=32'd186;
#400 value1=32'd264;value2=32'd280;
#400 value1=32'd299;value2=32'd314;
#400 value1=32'd320;value2=32'd321;
#400 value1=32'd326;value2=32'd331;
#400 value1=32'd332;value2=32'd335;
#400 value1=32'd336;value2=32'd466;
#400 value1=32'd494;value2=32'd530;
#400 value1=32'd127;value2=32'd187;
#400 value1=32'd265;value2=32'd290;
#400 value1=32'd307;value2=32'd314;
#400 value1=32'd320;value2=32'd322;
#400 value1=32'd327;value2=32'd330;
#400 value1=32'd333;value2=32'd337;
#400 value1=32'd338;value2=32'd467;
#400 value1=32'd495;value2=32'd531;
#400 value1=32'd128;value2=32'd188;
#400 value1=32'd266;value2=32'd280;
#400 value1=32'd299;value2=32'd323;
#400 value1=32'd325;value2=32'd328;
#400 value1=32'd330;value2=32'd333;
#400 value1=32'd339;value2=32'd468;
#400 value1=32'd496;value2=32'd532;
#400 value1=32'd129;value2=32'd189;
#400 value1=32'd267;value2=32'd290;
#400 value1=32'd307;value2=32'd324;
#400 value1=32'd325;value2=32'd329;
#400 value1=32'd331;value2=32'd332;
#400 value1=32'd339;value2=32'd469;
#400 value1=32'd497;value2=32'd533;
#400 value1=32'd190;value2=32'd268;
#400 value1=32'd282;value2=32'd291;
#400 value1=32'd301;value2=32'd308;
#400 value1=32'd315;value2=32'd316;
#400 value1=32'd321;value2=32'd322;
#400 value1=32'd336;value2=32'd337;
#400 value1=32'd470;value2=32'd498;
#400 value1=32'd534;value2=32'd550;
#400 value1=32'd191;value2=32'd269;
#400 value1=32'd281;value2=32'd283;
#400 value1=32'd300;value2=32'd302;
#400 value1=32'd317;value2=32'd323;
#400 value1=32'd326;value2=32'd330;
#400 value1=32'd336;value2=32'd337;
#400 value1=32'd471;value2=32'd499;
#400 value1=32'd535;value2=32'd551;
#400 value1=32'd192;value2=32'd270;
#400 value1=32'd284;value2=32'd291;
#400 value1=32'd303;value2=32'd308;
#400 value1=32'd318;value2=32'd324;
#400 value1=32'd326;value2=32'd330;
#400 value1=32'd334;value2=32'd335;
#400 value1=32'd338;value2=32'd339;
#400 value1=32'd472;value2=32'd500;
#400 value1=32'd536;value2=32'd552;
#400 value1=32'd193;value2=32'd271;
#400 value1=32'd282;value2=32'd293;
#400 value1=32'd301;value2=32'd310;
#400 value1=32'd317;value2=32'd323;
#400 value1=32'd327;value2=32'd331;
#400 value1=32'd334;value2=32'd335;
#400 value1=32'd338;value2=32'd339;
#400 value1=32'd473;value2=32'd501;
#400 value1=32'd537;value2=32'd553;
#400 value1=32'd194;value2=32'd272;
#400 value1=32'd292;value2=32'd294;
#400 value1=32'd309;value2=32'd311;
#400 value1=32'd318;value2=32'd324;
#400 value1=32'd327;value2=32'd331;
#400 value1=32'd336;value2=32'd337;
#400 value1=32'd474;value2=32'd502;
#400 value1=32'd538;value2=32'd554;
#400 value1=32'd195;value2=32'd273;
#400 value1=32'd284;value2=32'd293;
#400 value1=32'd303;value2=32'd310;
#400 value1=32'd328;value2=32'd329;
#400 value1=32'd332;value2=32'd333;
#400 value1=32'd336;value2=32'd337;
#400 value1=32'd475;value2=32'd503;
#400 value1=32'd539;value2=32'd555;
#400 value1=32'd40;value2=32'd50;
#400 value1=32'd131;value2=32'd141;
#400 value1=32'd208;value2=32'd274;
#400 value1=32'd341;value2=32'd346;
#400 value1=32'd348;value2=32'd350;
#400 value1=32'd356;value2=32'd358;
#400 value1=32'd400;value2=32'd402;
#400 value1=32'd41;value2=32'd51;
#400 value1=32'd132;value2=32'd142;
#400 value1=32'd208;value2=32'd274;
#400 value1=32'd340;value2=32'd347;
#400 value1=32'd349;value2=32'd364;
#400 value1=32'd366;value2=32'd395;
#400 value1=32'd408;value2=32'd410;
#400 value1=32'd39;value2=32'd42;
#400 value1=32'd52;value2=32'd133;
#400 value1=32'd143;value2=32'd208;
#400 value1=32'd343;value2=32'd344;
#400 value1=32'd346;value2=32'd347;
#400 value1=32'd359;value2=32'd371;
#400 value1=32'd373;value2=32'd396;
#400 value1=32'd415;value2=32'd417;
#400 value1=32'd43;value2=32'd53;
#400 value1=32'd130;value2=32'd134;
#400 value1=32'd144;value2=32'd274;
#400 value1=32'd342;value2=32'd345;
#400 value1=32'd346;value2=32'd347;
#400 value1=32'd360;value2=32'd377;
#400 value1=32'd379;value2=32'd397;
#400 value1=32'd421;value2=32'd423;
#400 value1=32'd39;value2=32'd44;
#400 value1=32'd54;value2=32'd135;
#400 value1=32'd145;value2=32'd208;
#400 value1=32'd342;value2=32'd345;
#400 value1=32'd348;value2=32'd349;
#400 value1=32'd361;value2=32'd382;
#400 value1=32'd384;value2=32'd398;
#400 value1=32'd426;value2=32'd428;
#400 value1=32'd45;value2=32'd55;
#400 value1=32'd130;value2=32'd136;
#400 value1=32'd146;value2=32'd274;
#400 value1=32'd343;value2=32'd344;
#400 value1=32'd348;value2=32'd349;
#400 value1=32'd362;value2=32'd386;
#400 value1=32'd388;value2=32'd399;
#400 value1=32'd430;value2=32'd432;
#400 value1=32'd46;value2=32'd56;
#400 value1=32'd137;value2=32'd147;
#400 value1=32'd340;value2=32'd342;
#400 value1=32'd343;value2=32'd347;
#400 value1=32'd348;value2=32'd363;
#400 value1=32'd389;value2=32'd391;
#400 value1=32'd400;value2=32'd435;
#400 value1=32'd47;value2=32'd57;
#400 value1=32'd138;value2=32'd148;
#400 value1=32'd341;value2=32'd342;
#400 value1=32'd343;value2=32'd346;
#400 value1=32'd349;value2=32'd364;
#400 value1=32'd393;value2=32'd401;
#400 value1=32'd434;value2=32'd437;
#400 value1=32'd48;value2=32'd58;
#400 value1=32'd139;value2=32'd149;
#400 value1=32'd340;value2=32'd344;
#400 value1=32'd345;value2=32'd346;
#400 value1=32'd349;value2=32'd365;
#400 value1=32'd392;value2=32'd394;
#400 value1=32'd402;value2=32'd435;
#400 value1=32'd49;value2=32'd59;
#400 value1=32'd140;value2=32'd150;
#400 value1=32'd341;value2=32'd344;
#400 value1=32'd345;value2=32'd347;
#400 value1=32'd348;value2=32'd366;
#400 value1=32'd393;value2=32'd403;
#400 value1=32'd436;value2=32'd439;
#400 value1=32'd60;value2=32'd151;
#400 value1=32'd209;value2=32'd210;
#400 value1=32'd275;value2=32'd276;
#400 value1=32'd340;value2=32'd356;
#400 value1=32'd358;value2=32'd363;
#400 value1=32'd365;value2=32'd395;
#400 value1=32'd444;value2=32'd446;
#400 value1=32'd40;value2=32'd61;
#400 value1=32'd152;value2=32'd209;
#400 value1=32'd211;value2=32'd277;
#400 value1=32'd352;value2=32'd353;
#400 value1=32'd355;value2=32'd356;
#400 value1=32'd359;value2=32'd370;
#400 value1=32'd372;value2=32'd396;
#400 value1=32'd451;value2=32'd453;
#400 value1=32'd62;value2=32'd131;
#400 value1=32'd153;value2=32'd212;
#400 value1=32'd275;value2=32'd278;
#400 value1=32'd351;value2=32'd354;
#400 value1=32'd355;value2=32'd356;
#400 value1=32'd360;value2=32'd376;
#400 value1=32'd378;value2=32'd397;
#400 value1=32'd457;value2=32'd459;
#400 value1=32'd40;value2=32'd63;
#400 value1=32'd154;value2=32'd209;
#400 value1=32'd213;value2=32'd279;
#400 value1=32'd351;value2=32'd354;
#400 value1=32'd357;value2=32'd358;
#400 value1=32'd361;value2=32'd381;
#400 value1=32'd383;value2=32'd398;
#400 value1=32'd462;value2=32'd464;
#400 value1=32'd64;value2=32'd131;
#400 value1=32'd155;value2=32'd214;
#400 value1=32'd275;value2=32'd280;
#400 value1=32'd352;value2=32'd353;
#400 value1=32'd357;value2=32'd358;
#400 value1=32'd362;value2=32'd385;
#400 value1=32'd387;value2=32'd399;
#400 value1=32'd466;value2=32'd468;
#400 value1=32'd65;value2=32'd156;
#400 value1=32'd215;value2=32'd281;
#400 value1=32'd351;value2=32'd352;
#400 value1=32'd356;value2=32'd357;
#400 value1=32'd363;value2=32'd390;
#400 value1=32'd400;value2=32'd471;
#400 value1=32'd66;value2=32'd157;
#400 value1=32'd216;value2=32'd282;
#400 value1=32'd340;value2=32'd350;
#400 value1=32'd351;value2=32'd352;
#400 value1=32'd355;value2=32'd358;
#400 value1=32'd364;value2=32'd389;
#400 value1=32'd392;value2=32'd401;
#400 value1=32'd470;value2=32'd473;
#400 value1=32'd67;value2=32'd158;
#400 value1=32'd217;value2=32'd283;
#400 value1=32'd353;value2=32'd354;
#400 value1=32'd355;value2=32'd358;
#400 value1=32'd365;value2=32'd390;
#400 value1=32'd402;value2=32'd471;
#400 value1=32'd68;value2=32'd159;
#400 value1=32'd218;value2=32'd284;
#400 value1=32'd340;value2=32'd350;
#400 value1=32'd353;value2=32'd354;
#400 value1=32'd356;value2=32'd357;
#400 value1=32'd366;value2=32'd391;
#400 value1=32'd394;value2=32'd403;
#400 value1=32'd472;value2=32'd475;
#400 value1=32'd41;value2=32'd69;
#400 value1=32'd160;value2=32'd210;
#400 value1=32'd211;value2=32'd277;
#400 value1=32'd342;value2=32'd351;
#400 value1=32'd360;value2=32'd361;
#400 value1=32'd363;value2=32'd364;
#400 value1=32'd371;value2=32'd373;
#400 value1=32'd404;value2=32'd440;
#400 value1=32'd479;value2=32'd481;
#400 value1=32'd70;value2=32'd132;
#400 value1=32'd161;value2=32'd212;
#400 value1=32'd276;value2=32'd278;
#400 value1=32'd343;value2=32'd352;
#400 value1=32'd359;value2=32'd362;
#400 value1=32'd363;value2=32'd364;
#400 value1=32'd377;value2=32'd379;
#400 value1=32'd405;value2=32'd441;
#400 value1=32'd485;value2=32'd487;
#400 value1=32'd41;value2=32'd71;
#400 value1=32'd162;value2=32'd210;
#400 value1=32'd213;value2=32'd279;
#400 value1=32'd344;value2=32'd353;
#400 value1=32'd359;value2=32'd362;
#400 value1=32'd365;value2=32'd366;
#400 value1=32'd382;value2=32'd384;
#400 value1=32'd406;value2=32'd442;
#400 value1=32'd490;value2=32'd492;
#400 value1=32'd72;value2=32'd132;
#400 value1=32'd163;value2=32'd214;
#400 value1=32'd276;value2=32'd280;
#400 value1=32'd345;value2=32'd354;
#400 value1=32'd360;value2=32'd361;
#400 value1=32'd365;value2=32'd366;
#400 value1=32'd386;value2=32'd388;
#400 value1=32'd407;value2=32'd443;
#400 value1=32'd494;value2=32'd496;
#400 value1=32'd73;value2=32'd164;
#400 value1=32'd215;value2=32'd281;
#400 value1=32'd346;value2=32'd350;
#400 value1=32'd355;value2=32'd359;
#400 value1=32'd360;value2=32'd364;
#400 value1=32'd365;value2=32'd389;
#400 value1=32'd391;value2=32'd408;
#400 value1=32'd444;value2=32'd499;
#400 value1=32'd74;value2=32'd165;
#400 value1=32'd216;value2=32'd282;
#400 value1=32'd341;value2=32'd347;
#400 value1=32'd356;value2=32'd359;
#400 value1=32'd360;value2=32'd363;
#400 value1=32'd366;value2=32'd393;
#400 value1=32'd409;value2=32'd445;
#400 value1=32'd498;value2=32'd501;
#400 value1=32'd75;value2=32'd166;
#400 value1=32'd217;value2=32'd283;
#400 value1=32'd348;value2=32'd350;
#400 value1=32'd357;value2=32'd361;
#400 value1=32'd362;value2=32'd363;
#400 value1=32'd366;value2=32'd392;
#400 value1=32'd394;value2=32'd410;
#400 value1=32'd446;value2=32'd499;
#400 value1=32'd76;value2=32'd167;
#400 value1=32'd218;value2=32'd284;
#400 value1=32'd341;value2=32'd349;
#400 value1=32'd358;value2=32'd361;
#400 value1=32'd362;value2=32'd364;
#400 value1=32'd365;value2=32'd393;
#400 value1=32'd411;value2=32'd447;
#400 value1=32'd500;value2=32'd503;
#400 value1=32'd43;value2=32'd77;
#400 value1=32'd133;value2=32'd168;
#400 value1=32'd212;value2=32'd277;
#400 value1=32'd369;value2=32'd370;
#400 value1=32'd371;value2=32'd374;
#400 value1=32'd376;value2=32'd377;
#400 value1=32'd412;value2=32'd448;
#400 value1=32'd506;value2=32'd508;
#400 value1=32'd42;value2=32'd44;
#400 value1=32'd78;value2=32'd169;
#400 value1=32'd211;value2=32'd213;
#400 value1=32'd369;value2=32'd372;
#400 value1=32'd373;value2=32'd374;
#400 value1=32'd381;value2=32'd382;
#400 value1=32'd413;value2=32'd449;
#400 value1=32'd511;value2=32'd513;
#400 value1=32'd45;value2=32'd79;
#400 value1=32'd133;value2=32'd170;
#400 value1=32'd214;value2=32'd277;
#400 value1=32'd367;value2=32'd368;
#400 value1=32'd372;value2=32'd373;
#400 value1=32'd375;value2=32'd380;
#400 value1=32'd385;value2=32'd386;
#400 value1=32'd414;value2=32'd450;
#400 value1=32'd515;value2=32'd517;
#400 value1=32'd46;value2=32'd80;
#400 value1=32'd171;value2=32'd215;
#400 value1=32'd351;value2=32'd367;
#400 value1=32'd371;value2=32'd372;
#400 value1=32'd376;value2=32'd381;
#400 value1=32'd389;value2=32'd415;
#400 value1=32'd451;value2=32'd520;
#400 value1=32'd47;value2=32'd81;
#400 value1=32'd172;value2=32'd216;
#400 value1=32'd342;value2=32'd359;
#400 value1=32'd367;value2=32'd370;
#400 value1=32'd373;value2=32'd377;
#400 value1=32'd382;value2=32'd389;
#400 value1=32'd416;value2=32'd452;
#400 value1=32'd519;value2=32'd522;
#400 value1=32'd48;value2=32'd82;
#400 value1=32'd173;value2=32'd217;
#400 value1=32'd351;value2=32'd368;
#400 value1=32'd369;value2=32'd370;
#400 value1=32'd373;value2=32'd378;
#400 value1=32'd383;value2=32'd390;
#400 value1=32'd392;value2=32'd417;
#400 value1=32'd453;value2=32'd520;
#400 value1=32'd49;value2=32'd83;
#400 value1=32'd174;value2=32'd218;
#400 value1=32'd342;value2=32'd359;
#400 value1=32'd368;value2=32'd369;
#400 value1=32'd371;value2=32'd372;
#400 value1=32'd379;value2=32'd384;
#400 value1=32'd391;value2=32'd393;
#400 value1=32'd418;value2=32'd454;
#400 value1=32'd521;value2=32'd524;
#400 value1=32'd43;value2=32'd84;
#400 value1=32'd135;value2=32'd175;
#400 value1=32'd212;value2=32'd279;
#400 value1=32'd367;value2=32'd368;
#400 value1=32'd375;value2=32'd378;
#400 value1=32'd379;value2=32'd380;
#400 value1=32'd381;value2=32'd382;
#400 value1=32'd419;value2=32'd455;
#400 value1=32'd526;value2=32'd528;
#400 value1=32'd85;value2=32'd134;
#400 value1=32'd136;value2=32'd176;
#400 value1=32'd278;value2=32'd280;
#400 value1=32'd369;value2=32'd374;
#400 value1=32'd378;value2=32'd379;
#400 value1=32'd385;value2=32'd386;
#400 value1=32'd420;value2=32'd456;
#400 value1=32'd530;value2=32'd532;
#400 value1=32'd86;value2=32'd137;
#400 value1=32'd177;value2=32'd281;
#400 value1=32'd352;value2=32'd367;
#400 value1=32'd370;value2=32'd377;
#400 value1=32'd378;value2=32'd385;
#400 value1=32'd389;value2=32'd421;
#400 value1=32'd457;value2=32'd535;
#400 value1=32'd87;value2=32'd138;
#400 value1=32'd178;value2=32'd282;
#400 value1=32'd343;value2=32'd360;
#400 value1=32'd367;value2=32'd371;
#400 value1=32'd376;value2=32'd379;
#400 value1=32'd386;value2=32'd389;
#400 value1=32'd422;value2=32'd458;
#400 value1=32'd534;value2=32'd537;
#400 value1=32'd88;value2=32'd139;
#400 value1=32'd179;value2=32'd283;
#400 value1=32'd352;value2=32'd372;
#400 value1=32'd374;value2=32'd375;
#400 value1=32'd376;value2=32'd379;
#400 value1=32'd387;value2=32'd390;
#400 value1=32'd392;value2=32'd423;
#400 value1=32'd459;value2=32'd535;
#400 value1=32'd89;value2=32'd140;
#400 value1=32'd180;value2=32'd284;
#400 value1=32'd343;value2=32'd360;
#400 value1=32'd373;value2=32'd374;
#400 value1=32'd375;value2=32'd377;
#400 value1=32'd378;value2=32'd388;
#400 value1=32'd391;value2=32'd393;
#400 value1=32'd424;value2=32'd460;
#400 value1=32'd536;value2=32'd539;
#400 value1=32'd45;value2=32'd90;
#400 value1=32'd135;value2=32'd181;
#400 value1=32'd214;value2=32'd279;
#400 value1=32'd369;value2=32'd374;
#400 value1=32'd383;value2=32'd384;
#400 value1=32'd387;value2=32'd388;
#400 value1=32'd425;value2=32'd461;
#400 value1=32'd540;value2=32'd542;
#400 value1=32'd46;value2=32'd91;
#400 value1=32'd182;value2=32'd215;
#400 value1=32'd353;value2=32'd368;
#400 value1=32'd370;value2=32'd374;
#400 value1=32'd382;value2=32'd383;
#400 value1=32'd385;value2=32'd390;
#400 value1=32'd391;value2=32'd426;
#400 value1=32'd462;value2=32'd545;
#400 value1=32'd47;value2=32'd92;
#400 value1=32'd183;value2=32'd216;
#400 value1=32'd344;value2=32'd361;
#400 value1=32'd368;value2=32'd371;
#400 value1=32'd374;value2=32'd381;
#400 value1=32'd384;value2=32'd386;
#400 value1=32'd392;value2=32'd393;
#400 value1=32'd427;value2=32'd463;
#400 value1=32'd544;value2=32'd547;
#400 value1=32'd48;value2=32'd93;
#400 value1=32'd184;value2=32'd217;
#400 value1=32'd353;value2=32'd372;
#400 value1=32'd380;value2=32'd381;
#400 value1=32'd384;value2=32'd387;
#400 value1=32'd394;value2=32'd428;
#400 value1=32'd464;value2=32'd545;
#400 value1=32'd49;value2=32'd94;
#400 value1=32'd185;value2=32'd218;
#400 value1=32'd344;value2=32'd361;
#400 value1=32'd373;value2=32'd380;
#400 value1=32'd382;value2=32'd383;
#400 value1=32'd388;value2=32'd394;
#400 value1=32'd429;value2=32'd465;
#400 value1=32'd546;value2=32'd549;
#400 value1=32'd95;value2=32'd137;
#400 value1=32'd186;value2=32'd281;
#400 value1=32'd354;value2=32'd369;
#400 value1=32'd375;value2=32'd376;
#400 value1=32'd381;value2=32'd386;
#400 value1=32'd387;value2=32'd390;
#400 value1=32'd391;value2=32'd430;
#400 value1=32'd466;value2=32'd551;
#400 value1=32'd96;value2=32'd138;
#400 value1=32'd187;value2=32'd282;
#400 value1=32'd345;value2=32'd362;
#400 value1=32'd369;value2=32'd375;
#400 value1=32'd377;value2=32'd382;
#400 value1=32'd385;value2=32'd388;
#400 value1=32'd392;value2=32'd393;
#400 value1=32'd431;value2=32'd467;
#400 value1=32'd550;value2=32'd553;
#400 value1=32'd97;value2=32'd139;
#400 value1=32'd188;value2=32'd283;
#400 value1=32'd354;value2=32'd378;
#400 value1=32'd380;value2=32'd383;
#400 value1=32'd385;value2=32'd388;
#400 value1=32'd394;value2=32'd432;
#400 value1=32'd468;value2=32'd551;
#400 value1=32'd98;value2=32'd140;
#400 value1=32'd189;value2=32'd284;
#400 value1=32'd345;value2=32'd362;
#400 value1=32'd379;value2=32'd380;
#400 value1=32'd384;value2=32'd386;
#400 value1=32'd387;value2=32'd394;
#400 value1=32'd433;value2=32'd469;
#400 value1=32'd552;value2=32'd555;
#400 value1=32'd99;value2=32'd190;
#400 value1=32'd346;value2=32'd356;
#400 value1=32'd363;value2=32'd370;
#400 value1=32'd371;value2=32'd376;
#400 value1=32'd377;value2=32'd391;
#400 value1=32'd392;value2=32'd434;
#400 value1=32'd470;value2=32'd556;
#400 value1=32'd100;value2=32'd191;
#400 value1=32'd355;value2=32'd357;
#400 value1=32'd372;value2=32'd378;
#400 value1=32'd381;value2=32'd385;
#400 value1=32'd391;value2=32'd392;
#400 value1=32'd435;value2=32'd471;
#400 value1=32'd101;value2=32'd192;
#400 value1=32'd346;value2=32'd358;
#400 value1=32'd363;value2=32'd373;
#400 value1=32'd379;value2=32'd381;
#400 value1=32'd385;value2=32'd389;
#400 value1=32'd390;value2=32'd393;
#400 value1=32'd394;value2=32'd436;
#400 value1=32'd472;value2=32'd558;
#400 value1=32'd102;value2=32'd193;
#400 value1=32'd348;value2=32'd356;
#400 value1=32'd365;value2=32'd372;
#400 value1=32'd378;value2=32'd382;
#400 value1=32'd386;value2=32'd389;
#400 value1=32'd390;value2=32'd393;
#400 value1=32'd394;value2=32'd437;
#400 value1=32'd473;value2=32'd556;
#400 value1=32'd103;value2=32'd194;
#400 value1=32'd347;value2=32'd349;
#400 value1=32'd364;value2=32'd366;
#400 value1=32'd373;value2=32'd379;
#400 value1=32'd382;value2=32'd386;
#400 value1=32'd391;value2=32'd392;
#400 value1=32'd438;value2=32'd474;
#400 value1=32'd557;value2=32'd559;
#400 value1=32'd104;value2=32'd195;
#400 value1=32'd348;value2=32'd358;
#400 value1=32'd365;value2=32'd383;
#400 value1=32'd384;value2=32'd387;
#400 value1=32'd388;value2=32'd391;
#400 value1=32'd392;value2=32'd439;
#400 value1=32'd475;value2=32'd558;
#400 value1=32'd60;value2=32'd151;
#400 value1=32'd219;value2=32'd220;
#400 value1=32'd285;value2=32'd286;
#400 value1=32'd341;value2=32'd350;
#400 value1=32'd401;value2=32'd403;
#400 value1=32'd408;value2=32'd410;
#400 value1=32'd445;value2=32'd447;
#400 value1=32'd50;value2=32'd61;
#400 value1=32'd152;value2=32'd219;
#400 value1=32'd221;value2=32'd287;
#400 value1=32'd342;value2=32'd351;
#400 value1=32'd397;value2=32'd398;
#400 value1=32'd400;value2=32'd401;
#400 value1=32'd404;value2=32'd415;
#400 value1=32'd417;value2=32'd440;
#400 value1=32'd452;value2=32'd454;
#400 value1=32'd62;value2=32'd141;
#400 value1=32'd153;value2=32'd222;
#400 value1=32'd285;value2=32'd288;
#400 value1=32'd343;value2=32'd352;
#400 value1=32'd396;value2=32'd399;
#400 value1=32'd400;value2=32'd401;
#400 value1=32'd405;value2=32'd421;
#400 value1=32'd423;value2=32'd441;
#400 value1=32'd458;value2=32'd460;
#400 value1=32'd50;value2=32'd63;
#400 value1=32'd154;value2=32'd219;
#400 value1=32'd223;value2=32'd289;
#400 value1=32'd344;value2=32'd353;
#400 value1=32'd396;value2=32'd399;
#400 value1=32'd402;value2=32'd403;
#400 value1=32'd406;value2=32'd426;
#400 value1=32'd428;value2=32'd442;
#400 value1=32'd463;value2=32'd465;
#400 value1=32'd64;value2=32'd141;
#400 value1=32'd155;value2=32'd224;
#400 value1=32'd285;value2=32'd290;
#400 value1=32'd345;value2=32'd354;
#400 value1=32'd397;value2=32'd398;
#400 value1=32'd402;value2=32'd403;
#400 value1=32'd407;value2=32'd430;
#400 value1=32'd432;value2=32'd443;
#400 value1=32'd467;value2=32'd469;
#400 value1=32'd65;value2=32'd156;
#400 value1=32'd225;value2=32'd291;
#400 value1=32'd340;value2=32'd346;
#400 value1=32'd355;value2=32'd396;
#400 value1=32'd397;value2=32'd401;
#400 value1=32'd402;value2=32'd408;
#400 value1=32'd435;value2=32'd444;
#400 value1=32'd470;value2=32'd472;
#400 value1=32'd66;value2=32'd157;
#400 value1=32'd226;value2=32'd292;
#400 value1=32'd347;value2=32'd356;
#400 value1=32'd395;value2=32'd396;
#400 value1=32'd397;value2=32'd400;
#400 value1=32'd403;value2=32'd409;
#400 value1=32'd434;value2=32'd437;
#400 value1=32'd445;value2=32'd474;
#400 value1=32'd67;value2=32'd158;
#400 value1=32'd227;value2=32'd293;
#400 value1=32'd340;value2=32'd348;
#400 value1=32'd357;value2=32'd398;
#400 value1=32'd399;value2=32'd400;
#400 value1=32'd403;value2=32'd410;
#400 value1=32'd435;value2=32'd446;
#400 value1=32'd473;value2=32'd475;
#400 value1=32'd68;value2=32'd159;
#400 value1=32'd228;value2=32'd294;
#400 value1=32'd349;value2=32'd358;
#400 value1=32'd395;value2=32'd398;
#400 value1=32'd399;value2=32'd401;
#400 value1=32'd402;value2=32'd411;
#400 value1=32'd436;value2=32'd439;
#400 value1=32'd447;value2=32'd474;
#400 value1=32'd51;value2=32'd69;
#400 value1=32'd160;value2=32'd220;
#400 value1=32'd221;value2=32'd287;
#400 value1=32'd359;value2=32'd396;
#400 value1=32'd405;value2=32'd406;
#400 value1=32'd408;value2=32'd409;
#400 value1=32'd416;value2=32'd418;
#400 value1=32'd480;value2=32'd482;
#400 value1=32'd70;value2=32'd142;
#400 value1=32'd161;value2=32'd222;
#400 value1=32'd286;value2=32'd288;
#400 value1=32'd360;value2=32'd397;
#400 value1=32'd404;value2=32'd407;
#400 value1=32'd408;value2=32'd409;
#400 value1=32'd422;value2=32'd424;
#400 value1=32'd486;value2=32'd488;
#400 value1=32'd51;value2=32'd71;
#400 value1=32'd162;value2=32'd220;
#400 value1=32'd223;value2=32'd289;
#400 value1=32'd361;value2=32'd398;
#400 value1=32'd404;value2=32'd407;
#400 value1=32'd410;value2=32'd411;
#400 value1=32'd427;value2=32'd429;
#400 value1=32'd491;value2=32'd493;
#400 value1=32'd72;value2=32'd142;
#400 value1=32'd163;value2=32'd224;
#400 value1=32'd286;value2=32'd290;
#400 value1=32'd362;value2=32'd399;
#400 value1=32'd405;value2=32'd406;
#400 value1=32'd410;value2=32'd411;
#400 value1=32'd431;value2=32'd433;
#400 value1=32'd495;value2=32'd497;
#400 value1=32'd73;value2=32'd164;
#400 value1=32'd225;value2=32'd291;
#400 value1=32'd341;value2=32'd363;
#400 value1=32'd395;value2=32'd400;
#400 value1=32'd404;value2=32'd405;
#400 value1=32'd409;value2=32'd410;
#400 value1=32'd434;value2=32'd436;
#400 value1=32'd498;value2=32'd500;
#400 value1=32'd74;value2=32'd165;
#400 value1=32'd226;value2=32'd292;
#400 value1=32'd364;value2=32'd401;
#400 value1=32'd404;value2=32'd405;
#400 value1=32'd408;value2=32'd411;
#400 value1=32'd438;value2=32'd502;
#400 value1=32'd75;value2=32'd166;
#400 value1=32'd227;value2=32'd293;
#400 value1=32'd341;value2=32'd365;
#400 value1=32'd395;value2=32'd402;
#400 value1=32'd406;value2=32'd407;
#400 value1=32'd408;value2=32'd411;
#400 value1=32'd437;value2=32'd439;
#400 value1=32'd501;value2=32'd503;
#400 value1=32'd76;value2=32'd167;
#400 value1=32'd228;value2=32'd294;
#400 value1=32'd366;value2=32'd403;
#400 value1=32'd406;value2=32'd407;
#400 value1=32'd409;value2=32'd410;
#400 value1=32'd438;value2=32'd502;
#400 value1=32'd53;value2=32'd77;
#400 value1=32'd143;value2=32'd168;
#400 value1=32'd222;value2=32'd287;
#400 value1=32'd367;value2=32'd414;
#400 value1=32'd415;value2=32'd416;
#400 value1=32'd419;value2=32'd421;
#400 value1=32'd422;value2=32'd476;
#400 value1=32'd507;value2=32'd509;
#400 value1=32'd52;value2=32'd54;
#400 value1=32'd78;value2=32'd169;
#400 value1=32'd221;value2=32'd223;
#400 value1=32'd368;value2=32'd414;
#400 value1=32'd417;value2=32'd418;
#400 value1=32'd419;value2=32'd426;
#400 value1=32'd427;value2=32'd477;
#400 value1=32'd512;value2=32'd514;
#400 value1=32'd55;value2=32'd79;
#400 value1=32'd143;value2=32'd170;
#400 value1=32'd224;value2=32'd287;
#400 value1=32'd369;value2=32'd412;
#400 value1=32'd413;value2=32'd417;
#400 value1=32'd418;value2=32'd420;
#400 value1=32'd425;value2=32'd430;
#400 value1=32'd431;value2=32'd478;
#400 value1=32'd516;value2=32'd518;
#400 value1=32'd56;value2=32'd80;
#400 value1=32'd171;value2=32'd225;
#400 value1=32'd342;value2=32'd370;
#400 value1=32'd396;value2=32'd412;
#400 value1=32'd416;value2=32'd417;
#400 value1=32'd421;value2=32'd426;
#400 value1=32'd434;value2=32'd479;
#400 value1=32'd519;value2=32'd521;
#400 value1=32'd57;value2=32'd81;
#400 value1=32'd172;value2=32'd226;
#400 value1=32'd371;value2=32'd404;
#400 value1=32'd412;value2=32'd415;
#400 value1=32'd418;value2=32'd422;
#400 value1=32'd427;value2=32'd434;
#400 value1=32'd480;value2=32'd523;
#400 value1=32'd58;value2=32'd82;
#400 value1=32'd173;value2=32'd227;
#400 value1=32'd342;value2=32'd372;
#400 value1=32'd396;value2=32'd413;
#400 value1=32'd414;value2=32'd415;
#400 value1=32'd418;value2=32'd423;
#400 value1=32'd428;value2=32'd435;
#400 value1=32'd437;value2=32'd481;
#400 value1=32'd522;value2=32'd524;
#400 value1=32'd59;value2=32'd83;
#400 value1=32'd174;value2=32'd228;
#400 value1=32'd373;value2=32'd404;
#400 value1=32'd413;value2=32'd414;
#400 value1=32'd416;value2=32'd417;
#400 value1=32'd424;value2=32'd429;
#400 value1=32'd436;value2=32'd438;
#400 value1=32'd482;value2=32'd523;
#400 value1=32'd53;value2=32'd84;
#400 value1=32'd145;value2=32'd175;
#400 value1=32'd222;value2=32'd289;
#400 value1=32'd374;value2=32'd412;
#400 value1=32'd413;value2=32'd420;
#400 value1=32'd423;value2=32'd424;
#400 value1=32'd425;value2=32'd426;
#400 value1=32'd427;value2=32'd483;
#400 value1=32'd527;value2=32'd529;
#400 value1=32'd85;value2=32'd144;
#400 value1=32'd146;value2=32'd176;
#400 value1=32'd288;value2=32'd290;
#400 value1=32'd375;value2=32'd414;
#400 value1=32'd419;value2=32'd423;
#400 value1=32'd424;value2=32'd430;
#400 value1=32'd431;value2=32'd484;
#400 value1=32'd531;value2=32'd533;
#400 value1=32'd86;value2=32'd147;
#400 value1=32'd177;value2=32'd291;
#400 value1=32'd343;value2=32'd376;
#400 value1=32'd397;value2=32'd412;
#400 value1=32'd415;value2=32'd422;
#400 value1=32'd423;value2=32'd430;
#400 value1=32'd434;value2=32'd485;
#400 value1=32'd534;value2=32'd536;
#400 value1=32'd87;value2=32'd148;
#400 value1=32'd178;value2=32'd292;
#400 value1=32'd377;value2=32'd405;
#400 value1=32'd412;value2=32'd416;
#400 value1=32'd421;value2=32'd424;
#400 value1=32'd431;value2=32'd434;
#400 value1=32'd486;value2=32'd538;
#400 value1=32'd88;value2=32'd149;
#400 value1=32'd179;value2=32'd293;
#400 value1=32'd343;value2=32'd378;
#400 value1=32'd397;value2=32'd417;
#400 value1=32'd419;value2=32'd420;
#400 value1=32'd421;value2=32'd424;
#400 value1=32'd432;value2=32'd435;
#400 value1=32'd437;value2=32'd487;
#400 value1=32'd537;value2=32'd539;
#400 value1=32'd89;value2=32'd150;
#400 value1=32'd180;value2=32'd294;
#400 value1=32'd379;value2=32'd405;
#400 value1=32'd418;value2=32'd419;
#400 value1=32'd420;value2=32'd422;
#400 value1=32'd423;value2=32'd433;
#400 value1=32'd436;value2=32'd438;
#400 value1=32'd488;value2=32'd538;
#400 value1=32'd55;value2=32'd90;
#400 value1=32'd145;value2=32'd181;
#400 value1=32'd224;value2=32'd289;
#400 value1=32'd380;value2=32'd414;
#400 value1=32'd419;value2=32'd428;
#400 value1=32'd429;value2=32'd432;
#400 value1=32'd433;value2=32'd489;
#400 value1=32'd541;value2=32'd543;
#400 value1=32'd56;value2=32'd91;
#400 value1=32'd182;value2=32'd225;
#400 value1=32'd344;value2=32'd381;
#400 value1=32'd398;value2=32'd413;
#400 value1=32'd415;value2=32'd419;
#400 value1=32'd427;value2=32'd428;
#400 value1=32'd430;value2=32'd435;
#400 value1=32'd436;value2=32'd490;
#400 value1=32'd544;value2=32'd546;
#400 value1=32'd57;value2=32'd92;
#400 value1=32'd183;value2=32'd226;
#400 value1=32'd382;value2=32'd406;
#400 value1=32'd413;value2=32'd416;
#400 value1=32'd419;value2=32'd426;
#400 value1=32'd429;value2=32'd431;
#400 value1=32'd437;value2=32'd438;
#400 value1=32'd491;value2=32'd548;
#400 value1=32'd58;value2=32'd93;
#400 value1=32'd184;value2=32'd227;
#400 value1=32'd344;value2=32'd383;
#400 value1=32'd398;value2=32'd417;
#400 value1=32'd425;value2=32'd426;
#400 value1=32'd429;value2=32'd432;
#400 value1=32'd439;value2=32'd492;
#400 value1=32'd547;value2=32'd549;
#400 value1=32'd59;value2=32'd94;
#400 value1=32'd185;value2=32'd228;
#400 value1=32'd384;value2=32'd406;
#400 value1=32'd418;value2=32'd425;
#400 value1=32'd427;value2=32'd428;
#400 value1=32'd433;value2=32'd439;
#400 value1=32'd493;value2=32'd548;
#400 value1=32'd95;value2=32'd147;
#400 value1=32'd186;value2=32'd291;
#400 value1=32'd345;value2=32'd385;
#400 value1=32'd399;value2=32'd414;
#400 value1=32'd420;value2=32'd421;
#400 value1=32'd426;value2=32'd431;
#400 value1=32'd432;value2=32'd435;
#400 value1=32'd436;value2=32'd494;
#400 value1=32'd550;value2=32'd552;
#400 value1=32'd96;value2=32'd148;
#400 value1=32'd187;value2=32'd292;
#400 value1=32'd386;value2=32'd407;
#400 value1=32'd414;value2=32'd420;
#400 value1=32'd422;value2=32'd427;
#400 value1=32'd430;value2=32'd433;
#400 value1=32'd437;value2=32'd438;
#400 value1=32'd495;value2=32'd554;
#400 value1=32'd97;value2=32'd149;
#400 value1=32'd188;value2=32'd293;
#400 value1=32'd345;value2=32'd387;
#400 value1=32'd399;value2=32'd423;
#400 value1=32'd425;value2=32'd428;
#400 value1=32'd430;value2=32'd433;
#400 value1=32'd439;value2=32'd496;
#400 value1=32'd553;value2=32'd555;
#400 value1=32'd98;value2=32'd150;
#400 value1=32'd189;value2=32'd294;
#400 value1=32'd388;value2=32'd407;
#400 value1=32'd424;value2=32'd425;
#400 value1=32'd429;value2=32'd431;
#400 value1=32'd432;value2=32'd439;
#400 value1=32'd497;value2=32'd554;
#400 value1=32'd99;value2=32'd190;
#400 value1=32'd347;value2=32'd389;
#400 value1=32'd401;value2=32'd408;
#400 value1=32'd415;value2=32'd416;
#400 value1=32'd421;value2=32'd422;
#400 value1=32'd436;value2=32'd437;
#400 value1=32'd498;value2=32'd557;
#400 value1=32'd100;value2=32'd191;
#400 value1=32'd346;value2=32'd348;
#400 value1=32'd390;value2=32'd400;
#400 value1=32'd402;value2=32'd417;
#400 value1=32'd423;value2=32'd426;
#400 value1=32'd430;value2=32'd436;
#400 value1=32'd437;value2=32'd499;
#400 value1=32'd556;value2=32'd558;
#400 value1=32'd101;value2=32'd192;
#400 value1=32'd349;value2=32'd391;
#400 value1=32'd403;value2=32'd408;
#400 value1=32'd418;value2=32'd424;
#400 value1=32'd426;value2=32'd430;
#400 value1=32'd434;value2=32'd435;
#400 value1=32'd438;value2=32'd439;
#400 value1=32'd500;value2=32'd557;
#400 value1=32'd102;value2=32'd193;
#400 value1=32'd347;value2=32'd392;
#400 value1=32'd401;value2=32'd410;
#400 value1=32'd417;value2=32'd423;
#400 value1=32'd427;value2=32'd431;
#400 value1=32'd434;value2=32'd435;
#400 value1=32'd438;value2=32'd439;
#400 value1=32'd501;value2=32'd559;
#400 value1=32'd103;value2=32'd194;
#400 value1=32'd393;value2=32'd409;
#400 value1=32'd411;value2=32'd418;
#400 value1=32'd424;value2=32'd427;
#400 value1=32'd431;value2=32'd436;
#400 value1=32'd437;value2=32'd502;
#400 value1=32'd104;value2=32'd195;
#400 value1=32'd349;value2=32'd394;
#400 value1=32'd403;value2=32'd410;
#400 value1=32'd428;value2=32'd429;
#400 value1=32'd432;value2=32'd433;
#400 value1=32'd436;value2=32'd437;
#400 value1=32'd503;value2=32'd559;
#400 value1=32'd60;value2=32'd229;
#400 value1=32'd230;value2=32'd238;
#400 value1=32'd296;value2=32'd304;
#400 value1=32'd359;value2=32'd396;
#400 value1=32'd441;value2=32'd442;
#400 value1=32'd444;value2=32'd445;
#400 value1=32'd452;value2=32'd454;
#400 value1=32'd479;value2=32'd481;
#400 value1=32'd151;value2=32'd231;
#400 value1=32'd239;value2=32'd295;
#400 value1=32'd297;value2=32'd305;
#400 value1=32'd360;value2=32'd397;
#400 value1=32'd440;value2=32'd443;
#400 value1=32'd444;value2=32'd445;
#400 value1=32'd458;value2=32'd460;
#400 value1=32'd485;value2=32'd487;
#400 value1=32'd60;value2=32'd229;
#400 value1=32'd232;value2=32'd240;
#400 value1=32'd298;value2=32'd306;
#400 value1=32'd361;value2=32'd398;
#400 value1=32'd440;value2=32'd443;
#400 value1=32'd446;value2=32'd447;
#400 value1=32'd463;value2=32'd465;
#400 value1=32'd490;value2=32'd492;
#400 value1=32'd151;value2=32'd233;
#400 value1=32'd241;value2=32'd295;
#400 value1=32'd299;value2=32'd307;
#400 value1=32'd362;value2=32'd399;
#400 value1=32'd441;value2=32'd442;
#400 value1=32'd446;value2=32'd447;
#400 value1=32'd467;value2=32'd469;
#400 value1=32'd494;value2=32'd496;
#400 value1=32'd234;value2=32'd242;
#400 value1=32'd300;value2=32'd308;
#400 value1=32'd350;value2=32'd363;
#400 value1=32'd400;value2=32'd440;
#400 value1=32'd441;value2=32'd445;
#400 value1=32'd446;value2=32'd470;
#400 value1=32'd472;value2=32'd499;
#400 value1=32'd235;value2=32'd243;
#400 value1=32'd301;value2=32'd309;
#400 value1=32'd364;value2=32'd395;
#400 value1=32'd401;value2=32'd440;
#400 value1=32'd441;value2=32'd444;
#400 value1=32'd447;value2=32'd474;
#400 value1=32'd498;value2=32'd501;
#400 value1=32'd236;value2=32'd244;
#400 value1=32'd302;value2=32'd310;
#400 value1=32'd350;value2=32'd365;
#400 value1=32'd402;value2=32'd442;
#400 value1=32'd443;value2=32'd444;
#400 value1=32'd447;value2=32'd473;
#400 value1=32'd475;value2=32'd499;
#400 value1=32'd237;value2=32'd245;
#400 value1=32'd303;value2=32'd311;
#400 value1=32'd366;value2=32'd395;
#400 value1=32'd403;value2=32'd442;
#400 value1=32'd443;value2=32'd445;
#400 value1=32'd446;value2=32'd474;
#400 value1=32'd500;value2=32'd503;
#400 value1=32'd62;value2=32'd152;
#400 value1=32'd231;value2=32'd246;
#400 value1=32'd296;value2=32'd312;
#400 value1=32'd367;value2=32'd450;
#400 value1=32'd451;value2=32'd452;
#400 value1=32'd455;value2=32'd457;
#400 value1=32'd458;value2=32'd476;
#400 value1=32'd506;value2=32'd508;
#400 value1=32'd61;value2=32'd63;
#400 value1=32'd230;value2=32'd232;
#400 value1=32'd247;value2=32'd313;
#400 value1=32'd368;value2=32'd450;
#400 value1=32'd453;value2=32'd454;
#400 value1=32'd455;value2=32'd462;
#400 value1=32'd463;value2=32'd477;
#400 value1=32'd511;value2=32'd513;
#400 value1=32'd64;value2=32'd152;
#400 value1=32'd233;value2=32'd248;
#400 value1=32'd296;value2=32'd314;
#400 value1=32'd369;value2=32'd448;
#400 value1=32'd449;value2=32'd453;
#400 value1=32'd454;value2=32'd456;
#400 value1=32'd461;value2=32'd466;
#400 value1=32'd467;value2=32'd478;
#400 value1=32'd515;value2=32'd517;
#400 value1=32'd65;value2=32'd234;
#400 value1=32'd249;value2=32'd315;
#400 value1=32'd351;value2=32'd370;
#400 value1=32'd448;value2=32'd452;
#400 value1=32'd453;value2=32'd457;
#400 value1=32'd462;value2=32'd470;
#400 value1=32'd479;value2=32'd520;
#400 value1=32'd66;value2=32'd235;
#400 value1=32'd250;value2=32'd316;
#400 value1=32'd371;value2=32'd396;
#400 value1=32'd440;value2=32'd448;
#400 value1=32'd451;value2=32'd454;
#400 value1=32'd458;value2=32'd463;
#400 value1=32'd470;value2=32'd480;
#400 value1=32'd519;value2=32'd522;
#400 value1=32'd67;value2=32'd236;
#400 value1=32'd251;value2=32'd317;
#400 value1=32'd351;value2=32'd372;
#400 value1=32'd449;value2=32'd450;
#400 value1=32'd451;value2=32'd454;
#400 value1=32'd459;value2=32'd464;
#400 value1=32'd471;value2=32'd473;
#400 value1=32'd481;value2=32'd520;
#400 value1=32'd68;value2=32'd237;
#400 value1=32'd252;value2=32'd318;
#400 value1=32'd373;value2=32'd396;
#400 value1=32'd440;value2=32'd449;
#400 value1=32'd450;value2=32'd452;
#400 value1=32'd453;value2=32'd460;
#400 value1=32'd465;value2=32'd472;
#400 value1=32'd474;value2=32'd482;
#400 value1=32'd521;value2=32'd524;
#400 value1=32'd62;value2=32'd154;
#400 value1=32'd231;value2=32'd253;
#400 value1=32'd298;value2=32'd319;
#400 value1=32'd374;value2=32'd448;
#400 value1=32'd449;value2=32'd456;
#400 value1=32'd459;value2=32'd460;
#400 value1=32'd461;value2=32'd462;
#400 value1=32'd463;value2=32'd483;
#400 value1=32'd526;value2=32'd528;
#400 value1=32'd153;value2=32'd155;
#400 value1=32'd254;value2=32'd297;
#400 value1=32'd299;value2=32'd320;
#400 value1=32'd375;value2=32'd450;
#400 value1=32'd455;value2=32'd459;
#400 value1=32'd460;value2=32'd466;
#400 value1=32'd467;value2=32'd484;
#400 value1=32'd530;value2=32'd532;
#400 value1=32'd156;value2=32'd255;
#400 value1=32'd300;value2=32'd321;
#400 value1=32'd352;value2=32'd376;
#400 value1=32'd448;value2=32'd451;
#400 value1=32'd458;value2=32'd459;
#400 value1=32'd466;value2=32'd470;
#400 value1=32'd485;value2=32'd535;
#400 value1=32'd157;value2=32'd256;
#400 value1=32'd301;value2=32'd322;
#400 value1=32'd377;value2=32'd397;
#400 value1=32'd441;value2=32'd448;
#400 value1=32'd452;value2=32'd457;
#400 value1=32'd460;value2=32'd467;
#400 value1=32'd470;value2=32'd486;
#400 value1=32'd534;value2=32'd537;
#400 value1=32'd158;value2=32'd257;
#400 value1=32'd302;value2=32'd323;
#400 value1=32'd352;value2=32'd378;
#400 value1=32'd453;value2=32'd455;
#400 value1=32'd456;value2=32'd457;
#400 value1=32'd460;value2=32'd468;
#400 value1=32'd471;value2=32'd473;
#400 value1=32'd487;value2=32'd535;
#400 value1=32'd159;value2=32'd258;
#400 value1=32'd303;value2=32'd324;
#400 value1=32'd379;value2=32'd397;
#400 value1=32'd441;value2=32'd454;
#400 value1=32'd455;value2=32'd456;
#400 value1=32'd458;value2=32'd459;
#400 value1=32'd469;value2=32'd472;
#400 value1=32'd474;value2=32'd488;
#400 value1=32'd536;value2=32'd539;
#400 value1=32'd64;value2=32'd154;
#400 value1=32'd233;value2=32'd259;
#400 value1=32'd298;value2=32'd325;
#400 value1=32'd380;value2=32'd450;
#400 value1=32'd455;value2=32'd464;
#400 value1=32'd465;value2=32'd468;
#400 value1=32'd469;value2=32'd489;
#400 value1=32'd540;value2=32'd542;
#400 value1=32'd65;value2=32'd234;
#400 value1=32'd260;value2=32'd326;
#400 value1=32'd353;value2=32'd381;
#400 value1=32'd449;value2=32'd451;
#400 value1=32'd455;value2=32'd463;
#400 value1=32'd464;value2=32'd466;
#400 value1=32'd471;value2=32'd472;
#400 value1=32'd490;value2=32'd545;
#400 value1=32'd66;value2=32'd235;
#400 value1=32'd261;value2=32'd327;
#400 value1=32'd382;value2=32'd398;
#400 value1=32'd442;value2=32'd449;
#400 value1=32'd452;value2=32'd455;
#400 value1=32'd462;value2=32'd465;
#400 value1=32'd467;value2=32'd473;
#400 value1=32'd474;value2=32'd491;
#400 value1=32'd544;value2=32'd547;
#400 value1=32'd67;value2=32'd236;
#400 value1=32'd262;value2=32'd328;
#400 value1=32'd353;value2=32'd383;
#400 value1=32'd453;value2=32'd461;
#400 value1=32'd462;value2=32'd465;
#400 value1=32'd468;value2=32'd475;
#400 value1=32'd492;value2=32'd545;
#400 value1=32'd68;value2=32'd237;
#400 value1=32'd263;value2=32'd329;
#400 value1=32'd384;value2=32'd398;
#400 value1=32'd442;value2=32'd454;
#400 value1=32'd461;value2=32'd463;
#400 value1=32'd464;value2=32'd469;
#400 value1=32'd475;value2=32'd493;
#400 value1=32'd546;value2=32'd549;
#400 value1=32'd156;value2=32'd264;
#400 value1=32'd300;value2=32'd330;
#400 value1=32'd354;value2=32'd385;
#400 value1=32'd450;value2=32'd456;
#400 value1=32'd457;value2=32'd462;
#400 value1=32'd467;value2=32'd468;
#400 value1=32'd471;value2=32'd472;
#400 value1=32'd494;value2=32'd551;
#400 value1=32'd157;value2=32'd265;
#400 value1=32'd301;value2=32'd331;
#400 value1=32'd386;value2=32'd399;
#400 value1=32'd443;value2=32'd450;
#400 value1=32'd456;value2=32'd458;
#400 value1=32'd463;value2=32'd466;
#400 value1=32'd469;value2=32'd473;
#400 value1=32'd474;value2=32'd495;
#400 value1=32'd550;value2=32'd553;
#400 value1=32'd158;value2=32'd266;
#400 value1=32'd302;value2=32'd332;
#400 value1=32'd354;value2=32'd387;
#400 value1=32'd459;value2=32'd461;
#400 value1=32'd464;value2=32'd466;
#400 value1=32'd469;value2=32'd475;
#400 value1=32'd496;value2=32'd551;
#400 value1=32'd159;value2=32'd267;
#400 value1=32'd303;value2=32'd333;
#400 value1=32'd388;value2=32'd399;
#400 value1=32'd443;value2=32'd460;
#400 value1=32'd461;value2=32'd465;
#400 value1=32'd467;value2=32'd468;
#400 value1=32'd475;value2=32'd497;
#400 value1=32'd552;value2=32'd555;
#400 value1=32'd268;value2=32'd334;
#400 value1=32'd356;value2=32'd389;
#400 value1=32'd400;value2=32'd444;
#400 value1=32'd451;value2=32'd452;
#400 value1=32'd457;value2=32'd458;
#400 value1=32'd472;value2=32'd473;
#400 value1=32'd498;value2=32'd556;
#400 value1=32'd269;value2=32'd335;
#400 value1=32'd355;value2=32'd357;
#400 value1=32'd390;value2=32'd453;
#400 value1=32'd459;value2=32'd462;
#400 value1=32'd466;value2=32'd472;
#400 value1=32'd473;value2=32'd499;
#400 value1=32'd270;value2=32'd336;
#400 value1=32'd358;value2=32'd391;
#400 value1=32'd400;value2=32'd444;
#400 value1=32'd454;value2=32'd460;
#400 value1=32'd462;value2=32'd466;
#400 value1=32'd470;value2=32'd471;
#400 value1=32'd474;value2=32'd475;
#400 value1=32'd500;value2=32'd558;
#400 value1=32'd271;value2=32'd337;
#400 value1=32'd356;value2=32'd392;
#400 value1=32'd402;value2=32'd446;
#400 value1=32'd453;value2=32'd459;
#400 value1=32'd463;value2=32'd467;
#400 value1=32'd470;value2=32'd471;
#400 value1=32'd474;value2=32'd475;
#400 value1=32'd501;value2=32'd556;
#400 value1=32'd272;value2=32'd338;
#400 value1=32'd393;value2=32'd401;
#400 value1=32'd403;value2=32'd445;
#400 value1=32'd447;value2=32'd454;
#400 value1=32'd460;value2=32'd463;
#400 value1=32'd467;value2=32'd472;
#400 value1=32'd473;value2=32'd502;
#400 value1=32'd557;value2=32'd559;
#400 value1=32'd273;value2=32'd339;
#400 value1=32'd358;value2=32'd394;
#400 value1=32'd402;value2=32'd446;
#400 value1=32'd464;value2=32'd465;
#400 value1=32'd468;value2=32'd469;
#400 value1=32'd472;value2=32'd473;
#400 value1=32'd503;value2=32'd558;
#400 value1=32'd70;value2=32'd160;
#400 value1=32'd239;value2=32'd246;
#400 value1=32'd304;value2=32'd312;
#400 value1=32'd412;value2=32'd448;
#400 value1=32'd478;value2=32'd479;
#400 value1=32'd480;value2=32'd483;
#400 value1=32'd485;value2=32'd486;
#400 value1=32'd507;value2=32'd509;
#400 value1=32'd69;value2=32'd71;
#400 value1=32'd238;value2=32'd240;
#400 value1=32'd247;value2=32'd313;
#400 value1=32'd413;value2=32'd449;
#400 value1=32'd478;value2=32'd481;
#400 value1=32'd482;value2=32'd483;
#400 value1=32'd490;value2=32'd491;
#400 value1=32'd512;value2=32'd514;
#400 value1=32'd72;value2=32'd160;
#400 value1=32'd241;value2=32'd248;
#400 value1=32'd304;value2=32'd314;
#400 value1=32'd414;value2=32'd450;
#400 value1=32'd476;value2=32'd477;
#400 value1=32'd481;value2=32'd482;
#400 value1=32'd484;value2=32'd489;
#400 value1=32'd494;value2=32'd495;
#400 value1=32'd516;value2=32'd518;
#400 value1=32'd73;value2=32'd242;
#400 value1=32'd249;value2=32'd315;
#400 value1=32'd359;value2=32'd415;
#400 value1=32'd440;value2=32'd451;
#400 value1=32'd476;value2=32'd480;
#400 value1=32'd481;value2=32'd485;
#400 value1=32'd490;value2=32'd498;
#400 value1=32'd519;value2=32'd521;
#400 value1=32'd74;value2=32'd243;
#400 value1=32'd250;value2=32'd316;
#400 value1=32'd404;value2=32'd416;
#400 value1=32'd452;value2=32'd476;
#400 value1=32'd479;value2=32'd482;
#400 value1=32'd486;value2=32'd491;
#400 value1=32'd498;value2=32'd523;
#400 value1=32'd75;value2=32'd244;
#400 value1=32'd251;value2=32'd317;
#400 value1=32'd359;value2=32'd417;
#400 value1=32'd440;value2=32'd453;
#400 value1=32'd477;value2=32'd478;
#400 value1=32'd479;value2=32'd482;
#400 value1=32'd487;value2=32'd492;
#400 value1=32'd499;value2=32'd501;
#400 value1=32'd522;value2=32'd524;
#400 value1=32'd76;value2=32'd245;
#400 value1=32'd252;value2=32'd318;
#400 value1=32'd404;value2=32'd418;
#400 value1=32'd454;value2=32'd477;
#400 value1=32'd478;value2=32'd480;
#400 value1=32'd481;value2=32'd488;
#400 value1=32'd493;value2=32'd500;
#400 value1=32'd502;value2=32'd523;
#400 value1=32'd70;value2=32'd162;
#400 value1=32'd239;value2=32'd253;
#400 value1=32'd306;value2=32'd319;
#400 value1=32'd419;value2=32'd455;
#400 value1=32'd476;value2=32'd477;
#400 value1=32'd484;value2=32'd487;
#400 value1=32'd488;value2=32'd489;
#400 value1=32'd490;value2=32'd491;
#400 value1=32'd527;value2=32'd529;
#400 value1=32'd161;value2=32'd163;
#400 value1=32'd254;value2=32'd305;
#400 value1=32'd307;value2=32'd320;
#400 value1=32'd420;value2=32'd456;
#400 value1=32'd478;value2=32'd483;
#400 value1=32'd487;value2=32'd488;
#400 value1=32'd494;value2=32'd495;
#400 value1=32'd531;value2=32'd533;
#400 value1=32'd164;value2=32'd255;
#400 value1=32'd308;value2=32'd321;
#400 value1=32'd360;value2=32'd421;
#400 value1=32'd441;value2=32'd457;
#400 value1=32'd476;value2=32'd479;
#400 value1=32'd486;value2=32'd487;
#400 value1=32'd494;value2=32'd498;
#400 value1=32'd534;value2=32'd536;
#400 value1=32'd165;value2=32'd256;
#400 value1=32'd309;value2=32'd322;
#400 value1=32'd405;value2=32'd422;
#400 value1=32'd458;value2=32'd476;
#400 value1=32'd480;value2=32'd485;
#400 value1=32'd488;value2=32'd495;
#400 value1=32'd498;value2=32'd538;
#400 value1=32'd166;value2=32'd257;
#400 value1=32'd310;value2=32'd323;
#400 value1=32'd360;value2=32'd423;
#400 value1=32'd441;value2=32'd459;
#400 value1=32'd481;value2=32'd483;
#400 value1=32'd484;value2=32'd485;
#400 value1=32'd488;value2=32'd496;
#400 value1=32'd499;value2=32'd501;
#400 value1=32'd537;value2=32'd539;
#400 value1=32'd167;value2=32'd258;
#400 value1=32'd311;value2=32'd324;
#400 value1=32'd405;value2=32'd424;
#400 value1=32'd460;value2=32'd482;
#400 value1=32'd483;value2=32'd484;
#400 value1=32'd486;value2=32'd487;
#400 value1=32'd497;value2=32'd500;
#400 value1=32'd502;value2=32'd538;
#400 value1=32'd72;value2=32'd162;
#400 value1=32'd241;value2=32'd259;
#400 value1=32'd306;value2=32'd325;
#400 value1=32'd425;value2=32'd461;
#400 value1=32'd478;value2=32'd483;
#400 value1=32'd492;value2=32'd493;
#400 value1=32'd496;value2=32'd497;
#400 value1=32'd541;value2=32'd543;
#400 value1=32'd73;value2=32'd242;
#400 value1=32'd260;value2=32'd326;
#400 value1=32'd361;value2=32'd426;
#400 value1=32'd442;value2=32'd462;
#400 value1=32'd477;value2=32'd479;
#400 value1=32'd483;value2=32'd491;
#400 value1=32'd492;value2=32'd494;
#400 value1=32'd499;value2=32'd500;
#400 value1=32'd544;value2=32'd546;
#400 value1=32'd74;value2=32'd243;
#400 value1=32'd261;value2=32'd327;
#400 value1=32'd406;value2=32'd427;
#400 value1=32'd463;value2=32'd477;
#400 value1=32'd480;value2=32'd483;
#400 value1=32'd490;value2=32'd493;
#400 value1=32'd495;value2=32'd501;
#400 value1=32'd502;value2=32'd548;
#400 value1=32'd75;value2=32'd244;
#400 value1=32'd262;value2=32'd328;
#400 value1=32'd361;value2=32'd428;
#400 value1=32'd442;value2=32'd464;
#400 value1=32'd481;value2=32'd489;
#400 value1=32'd490;value2=32'd493;
#400 value1=32'd496;value2=32'd503;
#400 value1=32'd547;value2=32'd549;
#400 value1=32'd76;value2=32'd245;
#400 value1=32'd263;value2=32'd329;
#400 value1=32'd406;value2=32'd429;
#400 value1=32'd465;value2=32'd482;
#400 value1=32'd489;value2=32'd491;
#400 value1=32'd492;value2=32'd497;
#400 value1=32'd503;value2=32'd548;
#400 value1=32'd164;value2=32'd264;
#400 value1=32'd308;value2=32'd330;
#400 value1=32'd362;value2=32'd430;
#400 value1=32'd443;value2=32'd466;
#400 value1=32'd478;value2=32'd484;
#400 value1=32'd485;value2=32'd490;
#400 value1=32'd495;value2=32'd496;
#400 value1=32'd499;value2=32'd500;
#400 value1=32'd550;value2=32'd552;
#400 value1=32'd165;value2=32'd265;
#400 value1=32'd309;value2=32'd331;
#400 value1=32'd407;value2=32'd431;
#400 value1=32'd467;value2=32'd478;
#400 value1=32'd484;value2=32'd486;
#400 value1=32'd491;value2=32'd494;
#400 value1=32'd497;value2=32'd501;
#400 value1=32'd502;value2=32'd554;
#400 value1=32'd166;value2=32'd266;
#400 value1=32'd310;value2=32'd332;
#400 value1=32'd362;value2=32'd432;
#400 value1=32'd443;value2=32'd468;
#400 value1=32'd487;value2=32'd489;
#400 value1=32'd492;value2=32'd494;
#400 value1=32'd497;value2=32'd503;
#400 value1=32'd553;value2=32'd555;
#400 value1=32'd167;value2=32'd267;
#400 value1=32'd311;value2=32'd333;
#400 value1=32'd407;value2=32'd433;
#400 value1=32'd469;value2=32'd488;
#400 value1=32'd489;value2=32'd493;
#400 value1=32'd495;value2=32'd496;
#400 value1=32'd503;value2=32'd554;
#400 value1=32'd268;value2=32'd334;
#400 value1=32'd364;value2=32'd408;
#400 value1=32'd434;value2=32'd445;
#400 value1=32'd470;value2=32'd479;
#400 value1=32'd480;value2=32'd485;
#400 value1=32'd486;value2=32'd500;
#400 value1=32'd501;value2=32'd557;
#400 value1=32'd269;value2=32'd335;
#400 value1=32'd363;value2=32'd365;
#400 value1=32'd435;value2=32'd444;
#400 value1=32'd446;value2=32'd471;
#400 value1=32'd481;value2=32'd487;
#400 value1=32'd490;value2=32'd494;
#400 value1=32'd500;value2=32'd501;
#400 value1=32'd556;value2=32'd558;
#400 value1=32'd270;value2=32'd336;
#400 value1=32'd366;value2=32'd408;
#400 value1=32'd436;value2=32'd447;
#400 value1=32'd472;value2=32'd482;
#400 value1=32'd488;value2=32'd490;
#400 value1=32'd494;value2=32'd498;
#400 value1=32'd499;value2=32'd502;
#400 value1=32'd503;value2=32'd557;
#400 value1=32'd271;value2=32'd337;
#400 value1=32'd364;value2=32'd410;
#400 value1=32'd437;value2=32'd445;
#400 value1=32'd473;value2=32'd481;
#400 value1=32'd487;value2=32'd491;
#400 value1=32'd495;value2=32'd498;
#400 value1=32'd499;value2=32'd502;
#400 value1=32'd503;value2=32'd559;
#400 value1=32'd272;value2=32'd338;
#400 value1=32'd409;value2=32'd411;
#400 value1=32'd438;value2=32'd474;
#400 value1=32'd482;value2=32'd488;
#400 value1=32'd491;value2=32'd495;
#400 value1=32'd500;value2=32'd501;
#400 value1=32'd273;value2=32'd339;
#400 value1=32'd366;value2=32'd410;
#400 value1=32'd439;value2=32'd447;
#400 value1=32'd475;value2=32'd492;
#400 value1=32'd493;value2=32'd496;
#400 value1=32'd497;value2=32'd500;
#400 value1=32'd501;value2=32'd559;
#400 value1=32'd77;value2=32'd84;
#400 value1=32'd169;value2=32'd246;
#400 value1=32'd253;value2=32'd313;
#400 value1=32'd505;value2=32'd508;
#400 value1=32'd509;value2=32'd510;
#400 value1=32'd511;value2=32'd512;
#400 value1=32'd526;value2=32'd527;
#400 value1=32'd85;value2=32'd168;
#400 value1=32'd170;value2=32'd254;
#400 value1=32'd312;value2=32'd314;
#400 value1=32'd504;value2=32'd508;
#400 value1=32'd509;value2=32'd515;
#400 value1=32'd516;value2=32'd525;
#400 value1=32'd530;value2=32'd531;
#400 value1=32'd86;value2=32'd171;
#400 value1=32'd255;value2=32'd315;
#400 value1=32'd367;value2=32'd448;
#400 value1=32'd507;value2=32'd508;
#400 value1=32'd515;value2=32'd519;
#400 value1=32'd526;value2=32'd534;
#400 value1=32'd87;value2=32'd172;
#400 value1=32'd256;value2=32'd316;
#400 value1=32'd412;value2=32'd476;
#400 value1=32'd506;value2=32'd509;
#400 value1=32'd516;value2=32'd519;
#400 value1=32'd527;value2=32'd534;
#400 value1=32'd88;value2=32'd173;
#400 value1=32'd257;value2=32'd317;
#400 value1=32'd367;value2=32'd448;
#400 value1=32'd504;value2=32'd505;
#400 value1=32'd506;value2=32'd509;
#400 value1=32'd517;value2=32'd520;
#400 value1=32'd522;value2=32'd528;
#400 value1=32'd535;value2=32'd537;
#400 value1=32'd89;value2=32'd174;
#400 value1=32'd258;value2=32'd318;
#400 value1=32'd412;value2=32'd476;
#400 value1=32'd504;value2=32'd505;
#400 value1=32'd507;value2=32'd508;
#400 value1=32'd518;value2=32'd521;
#400 value1=32'd523;value2=32'd529;
#400 value1=32'd536;value2=32'd538;
#400 value1=32'd79;value2=32'd90;
#400 value1=32'd169;value2=32'd248;
#400 value1=32'd259;value2=32'd313;
#400 value1=32'd504;value2=32'd513;
#400 value1=32'd514;value2=32'd517;
#400 value1=32'd518;value2=32'd525;
#400 value1=32'd540;value2=32'd541;
#400 value1=32'd80;value2=32'd91;
#400 value1=32'd249;value2=32'd260;
#400 value1=32'd368;value2=32'd449;
#400 value1=32'd504;value2=32'd512;
#400 value1=32'd513;value2=32'd515;
#400 value1=32'd520;value2=32'd521;
#400 value1=32'd526;value2=32'd544;
#400 value1=32'd81;value2=32'd92;
#400 value1=32'd250;value2=32'd261;
#400 value1=32'd413;value2=32'd477;
#400 value1=32'd504;value2=32'd511;
#400 value1=32'd514;value2=32'd516;
#400 value1=32'd522;value2=32'd523;
#400 value1=32'd527;value2=32'd544;
#400 value1=32'd82;value2=32'd93;
#400 value1=32'd251;value2=32'd262;
#400 value1=32'd368;value2=32'd449;
#400 value1=32'd510;value2=32'd511;
#400 value1=32'd514;value2=32'd517;
#400 value1=32'd524;value2=32'd528;
#400 value1=32'd545;value2=32'd547;
#400 value1=32'd83;value2=32'd94;
#400 value1=32'd252;value2=32'd263;
#400 value1=32'd413;value2=32'd477;
#400 value1=32'd510;value2=32'd512;
#400 value1=32'd513;value2=32'd518;
#400 value1=32'd524;value2=32'd529;
#400 value1=32'd546;value2=32'd548;
#400 value1=32'd95;value2=32'd171;
#400 value1=32'd264;value2=32'd315;
#400 value1=32'd369;value2=32'd450;
#400 value1=32'd505;value2=32'd506;
#400 value1=32'd511;value2=32'd516;
#400 value1=32'd517;value2=32'd520;
#400 value1=32'd521;value2=32'd530;
#400 value1=32'd540;value2=32'd550;
#400 value1=32'd96;value2=32'd172;
#400 value1=32'd265;value2=32'd316;
#400 value1=32'd414;value2=32'd478;
#400 value1=32'd505;value2=32'd507;
#400 value1=32'd512;value2=32'd515;
#400 value1=32'd518;value2=32'd522;
#400 value1=32'd523;value2=32'd531;
#400 value1=32'd541;value2=32'd550;
#400 value1=32'd97;value2=32'd173;
#400 value1=32'd266;value2=32'd317;
#400 value1=32'd369;value2=32'd450;
#400 value1=32'd508;value2=32'd510;
#400 value1=32'd513;value2=32'd515;
#400 value1=32'd518;value2=32'd524;
#400 value1=32'd532;value2=32'd542;
#400 value1=32'd551;value2=32'd553;
#400 value1=32'd98;value2=32'd174;
#400 value1=32'd267;value2=32'd318;
#400 value1=32'd414;value2=32'd478;
#400 value1=32'd509;value2=32'd510;
#400 value1=32'd514;value2=32'd516;
#400 value1=32'd517;value2=32'd524;
#400 value1=32'd533;value2=32'd543;
#400 value1=32'd552;value2=32'd554;
#400 value1=32'd99;value2=32'd268;
#400 value1=32'd371;value2=32'd415;
#400 value1=32'd452;value2=32'd479;
#400 value1=32'd506;value2=32'd507;
#400 value1=32'd521;value2=32'd522;
#400 value1=32'd534;value2=32'd544;
#400 value1=32'd100;value2=32'd269;
#400 value1=32'd370;value2=32'd372;
#400 value1=32'd451;value2=32'd453;
#400 value1=32'd508;value2=32'd511;
#400 value1=32'd515;value2=32'd521;
#400 value1=32'd522;value2=32'd535;
#400 value1=32'd545;value2=32'd556;
#400 value1=32'd101;value2=32'd270;
#400 value1=32'd373;value2=32'd415;
#400 value1=32'd454;value2=32'd479;
#400 value1=32'd509;value2=32'd511;
#400 value1=32'd515;value2=32'd519;
#400 value1=32'd520;value2=32'd523;
#400 value1=32'd524;value2=32'd536;
#400 value1=32'd546;value2=32'd557;
#400 value1=32'd102;value2=32'd271;
#400 value1=32'd371;value2=32'd417;
#400 value1=32'd452;value2=32'd481;
#400 value1=32'd508;value2=32'd512;
#400 value1=32'd516;value2=32'd519;
#400 value1=32'd520;value2=32'd523;
#400 value1=32'd524;value2=32'd537;
#400 value1=32'd547;value2=32'd556;
#400 value1=32'd103;value2=32'd272;
#400 value1=32'd416;value2=32'd418;
#400 value1=32'd480;value2=32'd482;
#400 value1=32'd509;value2=32'd512;
#400 value1=32'd516;value2=32'd521;
#400 value1=32'd522;value2=32'd538;
#400 value1=32'd548;value2=32'd557;
#400 value1=32'd104;value2=32'd273;
#400 value1=32'd373;value2=32'd417;
#400 value1=32'd454;value2=32'd481;
#400 value1=32'd513;value2=32'd514;
#400 value1=32'd517;value2=32'd518;
#400 value1=32'd521;value2=32'd522;
#400 value1=32'd539;value2=32'd549;
#400 value1=32'd558;value2=32'd559;
#400 value1=32'd85;value2=32'd175;
#400 value1=32'd181;value2=32'd254;
#400 value1=32'd319;value2=32'd325;
#400 value1=32'd505;value2=32'd510;
#400 value1=32'd528;value2=32'd529;
#400 value1=32'd532;value2=32'd533;
#400 value1=32'd540;value2=32'd541;
#400 value1=32'd86;value2=32'd182;
#400 value1=32'd255;value2=32'd326;
#400 value1=32'd374;value2=32'd455;
#400 value1=32'd504;value2=32'd506;
#400 value1=32'd511;value2=32'd527;
#400 value1=32'd528;value2=32'd530;
#400 value1=32'd535;value2=32'd536;
#400 value1=32'd540;value2=32'd544;
#400 value1=32'd87;value2=32'd183;
#400 value1=32'd256;value2=32'd327;
#400 value1=32'd419;value2=32'd483;
#400 value1=32'd504;value2=32'd507;
#400 value1=32'd512;value2=32'd526;
#400 value1=32'd529;value2=32'd531;
#400 value1=32'd537;value2=32'd538;
#400 value1=32'd541;value2=32'd544;
#400 value1=32'd88;value2=32'd184;
#400 value1=32'd257;value2=32'd328;
#400 value1=32'd374;value2=32'd455;
#400 value1=32'd508;value2=32'd513;
#400 value1=32'd525;value2=32'd526;
#400 value1=32'd529;value2=32'd532;
#400 value1=32'd539;value2=32'd542;
#400 value1=32'd545;value2=32'd547;
#400 value1=32'd89;value2=32'd185;
#400 value1=32'd258;value2=32'd329;
#400 value1=32'd419;value2=32'd483;
#400 value1=32'd509;value2=32'd514;
#400 value1=32'd525;value2=32'd527;
#400 value1=32'd528;value2=32'd533;
#400 value1=32'd539;value2=32'd543;
#400 value1=32'd546;value2=32'd548;
#400 value1=32'd177;value2=32'd186;
#400 value1=32'd321;value2=32'd330;
#400 value1=32'd375;value2=32'd456;
#400 value1=32'd505;value2=32'd515;
#400 value1=32'd526;value2=32'd531;
#400 value1=32'd532;value2=32'd535;
#400 value1=32'd536;value2=32'd550;
#400 value1=32'd178;value2=32'd187;
#400 value1=32'd322;value2=32'd331;
#400 value1=32'd420;value2=32'd484;
#400 value1=32'd505;value2=32'd516;
#400 value1=32'd527;value2=32'd530;
#400 value1=32'd533;value2=32'd537;
#400 value1=32'd538;value2=32'd550;
#400 value1=32'd179;value2=32'd188;
#400 value1=32'd323;value2=32'd332;
#400 value1=32'd375;value2=32'd456;
#400 value1=32'd517;value2=32'd525;
#400 value1=32'd528;value2=32'd530;
#400 value1=32'd533;value2=32'd539;
#400 value1=32'd551;value2=32'd553;
#400 value1=32'd180;value2=32'd189;
#400 value1=32'd324;value2=32'd333;
#400 value1=32'd420;value2=32'd484;
#400 value1=32'd518;value2=32'd525;
#400 value1=32'd529;value2=32'd531;
#400 value1=32'd532;value2=32'd539;
#400 value1=32'd552;value2=32'd554;
#400 value1=32'd190;value2=32'd334;
#400 value1=32'd377;value2=32'd421;
#400 value1=32'd458;value2=32'd485;
#400 value1=32'd506;value2=32'd507;
#400 value1=32'd519;value2=32'd536;
#400 value1=32'd537;value2=32'd550;
#400 value1=32'd191;value2=32'd335;
#400 value1=32'd376;value2=32'd378;
#400 value1=32'd457;value2=32'd459;
#400 value1=32'd508;value2=32'd520;
#400 value1=32'd526;value2=32'd530;
#400 value1=32'd536;value2=32'd537;
#400 value1=32'd551;value2=32'd556;
#400 value1=32'd192;value2=32'd336;
#400 value1=32'd379;value2=32'd421;
#400 value1=32'd460;value2=32'd485;
#400 value1=32'd509;value2=32'd521;
#400 value1=32'd526;value2=32'd530;
#400 value1=32'd534;value2=32'd535;
#400 value1=32'd538;value2=32'd539;
#400 value1=32'd552;value2=32'd557;
#400 value1=32'd193;value2=32'd337;
#400 value1=32'd377;value2=32'd423;
#400 value1=32'd458;value2=32'd487;
#400 value1=32'd508;value2=32'd522;
#400 value1=32'd527;value2=32'd531;
#400 value1=32'd534;value2=32'd535;
#400 value1=32'd538;value2=32'd539;
#400 value1=32'd553;value2=32'd556;
#400 value1=32'd194;value2=32'd338;
#400 value1=32'd422;value2=32'd424;
#400 value1=32'd486;value2=32'd488;
#400 value1=32'd509;value2=32'd523;
#400 value1=32'd527;value2=32'd531;
#400 value1=32'd536;value2=32'd537;
#400 value1=32'd554;value2=32'd557;
#400 value1=32'd195;value2=32'd339;
#400 value1=32'd379;value2=32'd423;
#400 value1=32'd460;value2=32'd487;
#400 value1=32'd524;value2=32'd528;
#400 value1=32'd529;value2=32'd532;
#400 value1=32'd533;value2=32'd536;
#400 value1=32'd537;value2=32'd555;
#400 value1=32'd558;value2=32'd559;
#400 value1=32'd95;value2=32'd182;
#400 value1=32'd264;value2=32'd326;
#400 value1=32'd380;value2=32'd461;
#400 value1=32'd510;value2=32'd515;
#400 value1=32'd525;value2=32'd526;
#400 value1=32'd541;value2=32'd542;
#400 value1=32'd545;value2=32'd546;
#400 value1=32'd551;value2=32'd552;
#400 value1=32'd96;value2=32'd183;
#400 value1=32'd265;value2=32'd327;
#400 value1=32'd425;value2=32'd489;
#400 value1=32'd510;value2=32'd516;
#400 value1=32'd525;value2=32'd527;
#400 value1=32'd540;value2=32'd543;
#400 value1=32'd547;value2=32'd548;
#400 value1=32'd553;value2=32'd554;
#400 value1=32'd97;value2=32'd184;
#400 value1=32'd266;value2=32'd328;
#400 value1=32'd380;value2=32'd461;
#400 value1=32'd517;value2=32'd528;
#400 value1=32'd540;value2=32'd543;
#400 value1=32'd549;value2=32'd555;
#400 value1=32'd98;value2=32'd185;
#400 value1=32'd267;value2=32'd329;
#400 value1=32'd425;value2=32'd489;
#400 value1=32'd518;value2=32'd529;
#400 value1=32'd541;value2=32'd542;
#400 value1=32'd549;value2=32'd555;
#400 value1=32'd99;value2=32'd268;
#400 value1=32'd382;value2=32'd426;
#400 value1=32'd463;value2=32'd490;
#400 value1=32'd511;value2=32'd512;
#400 value1=32'd519;value2=32'd526;
#400 value1=32'd527;value2=32'd546;
#400 value1=32'd547;value2=32'd550;
#400 value1=32'd556;value2=32'd557;
#400 value1=32'd100;value2=32'd269;
#400 value1=32'd381;value2=32'd383;
#400 value1=32'd462;value2=32'd464;
#400 value1=32'd513;value2=32'd520;
#400 value1=32'd528;value2=32'd540;
#400 value1=32'd546;value2=32'd547;
#400 value1=32'd551;value2=32'd558;
#400 value1=32'd101;value2=32'd270;
#400 value1=32'd384;value2=32'd426;
#400 value1=32'd465;value2=32'd490;
#400 value1=32'd514;value2=32'd521;
#400 value1=32'd529;value2=32'd540;
#400 value1=32'd544;value2=32'd545;
#400 value1=32'd548;value2=32'd549;
#400 value1=32'd552;value2=32'd558;
#400 value1=32'd102;value2=32'd271;
#400 value1=32'd382;value2=32'd428;
#400 value1=32'd463;value2=32'd492;
#400 value1=32'd513;value2=32'd522;
#400 value1=32'd528;value2=32'd541;
#400 value1=32'd544;value2=32'd545;
#400 value1=32'd548;value2=32'd549;
#400 value1=32'd553;value2=32'd559;
#400 value1=32'd103;value2=32'd272;
#400 value1=32'd427;value2=32'd429;
#400 value1=32'd491;value2=32'd493;
#400 value1=32'd514;value2=32'd523;
#400 value1=32'd529;value2=32'd541;
#400 value1=32'd546;value2=32'd547;
#400 value1=32'd554;value2=32'd559;
#400 value1=32'd104;value2=32'd273;
#400 value1=32'd384;value2=32'd428;
#400 value1=32'd465;value2=32'd492;
#400 value1=32'd524;value2=32'd542;
#400 value1=32'd543;value2=32'd546;
#400 value1=32'd547;value2=32'd555;
#400 value1=32'd190;value2=32'd334;
#400 value1=32'd386;value2=32'd430;
#400 value1=32'd467;value2=32'd494;
#400 value1=32'd515;value2=32'd516;
#400 value1=32'd530;value2=32'd531;
#400 value1=32'd534;value2=32'd544;
#400 value1=32'd552;value2=32'd553;
#400 value1=32'd556;value2=32'd557;
#400 value1=32'd191;value2=32'd335;
#400 value1=32'd385;value2=32'd387;
#400 value1=32'd466;value2=32'd468;
#400 value1=32'd517;value2=32'd532;
#400 value1=32'd535;value2=32'd540;
#400 value1=32'd545;value2=32'd552;
#400 value1=32'd553;value2=32'd558;
#400 value1=32'd192;value2=32'd336;
#400 value1=32'd388;value2=32'd430;
#400 value1=32'd469;value2=32'd494;
#400 value1=32'd518;value2=32'd533;
#400 value1=32'd536;value2=32'd540;
#400 value1=32'd546;value2=32'd550;
#400 value1=32'd551;value2=32'd554;
#400 value1=32'd555;value2=32'd558;
#400 value1=32'd193;value2=32'd337;
#400 value1=32'd386;value2=32'd432;
#400 value1=32'd467;value2=32'd496;
#400 value1=32'd517;value2=32'd532;
#400 value1=32'd537;value2=32'd541;
#400 value1=32'd547;value2=32'd550;
#400 value1=32'd551;value2=32'd554;
#400 value1=32'd555;value2=32'd559;
#400 value1=32'd194;value2=32'd338;
#400 value1=32'd431;value2=32'd433;
#400 value1=32'd495;value2=32'd497;
#400 value1=32'd518;value2=32'd533;
#400 value1=32'd538;value2=32'd541;
#400 value1=32'd548;value2=32'd552;
#400 value1=32'd553;value2=32'd559;
#400 value1=32'd195;value2=32'd339;
#400 value1=32'd388;value2=32'd432;
#400 value1=32'd469;value2=32'd496;
#400 value1=32'd539;value2=32'd542;
#400 value1=32'd543;value2=32'd549;
#400 value1=32'd552;value2=32'd553;
#400 value1=32'd389;value2=32'd392;
#400 value1=32'd435;value2=32'd470;
#400 value1=32'd473;value2=32'd499;
#400 value1=32'd520;value2=32'd522;
#400 value1=32'd535;value2=32'd537;
#400 value1=32'd544;value2=32'd550;
#400 value1=32'd557;value2=32'd558;
#400 value1=32'd393;value2=32'd434;
#400 value1=32'd436;value2=32'd474;
#400 value1=32'd498;value2=32'd500;
#400 value1=32'd521;value2=32'd523;
#400 value1=32'd536;value2=32'd538;
#400 value1=32'd544;value2=32'd550;
#400 value1=32'd556;value2=32'd559;
#400 value1=32'd391;value2=32'd394;
#400 value1=32'd435;value2=32'd472;
#400 value1=32'd475;value2=32'd499;
#400 value1=32'd524;value2=32'd539;
#400 value1=32'd545;value2=32'd546;
#400 value1=32'd551;value2=32'd552;
#400 value1=32'd556;value2=32'd559;
#400 value1=32'd393;value2=32'd437;
#400 value1=32'd439;value2=32'd474;
#400 value1=32'd501;value2=32'd503;
#400 value1=32'd524;value2=32'd539;
#400 value1=32'd547;value2=32'd548;
#400 value1=32'd553;value2=32'd554;
#400 value1=32'd557;value2=32'd558;
//rowpointer
#400 value1=32'd0;value2=32'd14;
#400 value1=32'd28;value2=32'd40;
#400 value1=32'd52;value2=32'd68;
#400 value1=32'd84;value2=32'd98;
#400 value1=32'd112;value2=32'd126;
#400 value1=32'd140;value2=32'd156;
#400 value1=32'd172;value2=32'd188;
#400 value1=32'd204;value2=32'd218;
#400 value1=32'd232;value2=32'd246;
#400 value1=32'd260;value2=32'd274;
#400 value1=32'd286;value2=32'd302;
#400 value1=32'd314;value2=32'd330;
#400 value1=32'd346;value2=32'd362;
#400 value1=32'd378;value2=32'd394;
#400 value1=32'd410;value2=32'd426;
#400 value1=32'd442;value2=32'd458;
#400 value1=32'd474;value2=32'd490;
#400 value1=32'd506;value2=32'd522;
#400 value1=32'd540;value2=32'd558;
#400 value1=32'd576;value2=32'd594;
#400 value1=32'd606;value2=32'd620;
#400 value1=32'd636;value2=32'd650;
#400 value1=32'd666;value2=32'd680;
#400 value1=32'd696;value2=32'd710;
#400 value1=32'd726;value2=32'd740;
#400 value1=32'd756;value2=32'd772;
#400 value1=32'd786;value2=32'd800;
#400 value1=32'd816;value2=32'd830;
#400 value1=32'd846;value2=32'd862;
#400 value1=32'd876;value2=32'd892;
#400 value1=32'd906;value2=32'd922;
#400 value1=32'd938;value2=32'd956;
#400 value1=32'd972;value2=32'd990;
#400 value1=32'd1006;value2=32'd1024;
#400 value1=32'd1040;value2=32'd1058;
#400 value1=32'd1074;value2=32'd1092;
#400 value1=32'd1108;value2=32'd1126;
#400 value1=32'd1144;value2=32'd1160;
#400 value1=32'd1178;value2=32'd1194;
#400 value1=32'd1208;value2=32'd1220;
#400 value1=32'd1236;value2=32'd1250;
#400 value1=32'd1264;value2=32'd1280;
#400 value1=32'd1296;value2=32'd1312;
#400 value1=32'd1328;value2=32'd1344;
#400 value1=32'd1360;value2=32'd1378;
#400 value1=32'd1396;value2=32'd1410;
#400 value1=32'd1426;value2=32'd1442;
#400 value1=32'd1456;value2=32'd1470;
#400 value1=32'd1488;value2=32'd1506;
#400 value1=32'd1522;value2=32'd1538;
#400 value1=32'd1554;value2=32'd1570;
#400 value1=32'd1588;value2=32'd1606;
#400 value1=32'd1622;value2=32'd1638;
#400 value1=32'd1652;value2=32'd1668;
#400 value1=32'd1684;value2=32'd1700;
#400 value1=32'd1716;value2=32'd1732;
#400 value1=32'd1748;value2=32'd1764;
#400 value1=32'd1780;value2=32'd1798;
#400 value1=32'd1816;value2=32'd1834;
#400 value1=32'd1852;value2=32'd1866;
#400 value1=32'd1880;value2=32'd1894;
#400 value1=32'd1908;value2=32'd1924;
#400 value1=32'd1936;value2=32'd1952;
#400 value1=32'd1964;value2=32'd1980;
#400 value1=32'd1996;value2=32'd2012;
#400 value1=32'd2028;value2=32'd2040;
#400 value1=32'd2054;value2=32'd2070;
#400 value1=32'd2086;value2=32'd2100;
#400 value1=32'd2116;value2=32'd2130;
#400 value1=32'd2144;value2=32'd2160;
#400 value1=32'd2174;value2=32'd2190;
#400 value1=32'd2206;value2=32'd2220;
#400 value1=32'd2236;value2=32'd2250;
#400 value1=32'd2266;value2=32'd2280;
#400 value1=32'd2296;value2=32'd2310;
#400 value1=32'd2326;value2=32'd2340;
#400 value1=32'd2356;value2=32'd2374;
#400 value1=32'd2390;value2=32'd2408;
#400 value1=32'd2424;value2=32'd2440;
#400 value1=32'd2458;value2=32'd2474;
#400 value1=32'd2492;value2=32'd2510;
#400 value1=32'd2526;value2=32'd2544;
#400 value1=32'd2560;value2=32'd2578;
#400 value1=32'd2594;value2=32'd2612;
#400 value1=32'd2628;value2=32'd2642;
#400 value1=32'd2658;value2=32'd2674;
#400 value1=32'd2690;value2=32'd2706;
#400 value1=32'd2724;value2=32'd2742;
#400 value1=32'd2758;value2=32'd2770;
#400 value1=32'd2784;value2=32'd2798;
#400 value1=32'd2814;value2=32'd2830;
#400 value1=32'd2844;value2=32'd2862;
#400 value1=32'd2880;value2=32'd2896;
#400 value1=32'd2912;value2=32'd2928;
#400 value1=32'd2944;value2=32'd2958;
#400 value1=32'd2972;value2=32'd2988;
#400 value1=32'd3004;value2=32'd3022;
#400 value1=32'd3040;value2=32'd3056;
#400 value1=32'd3072;value2=32'd3088;
#400 value1=32'd3104;value2=32'd3116;
#400 value1=32'd3128;value2=32'd3142;
#400 value1=32'd3156;value2=32'd3170;
#400 value1=32'd3184;value2=32'd3200;
#400 value1=32'd3216;value2=32'd3232;
#400 value1=32'd3248;value2=32'd3264;
#400 value1=32'd3278;value2=32'd3294;
#400 value1=32'd3310;value2=32'd3328;
#400 value1=32'd3344;value2=32'd3362;
#400 value1=32'd3378;value2=32'd3396;
#400 value1=32'd3412;value2=32'd3430;
#400 value1=32'd3446;value2=32'd3460;
#400 value1=32'd3476;value2=32'd3494;
#400 value1=32'd3510;value2=32'd3528;
#400 value1=32'd3546;value2=32'd3562;
#400 value1=32'd3580;value2=32'd3596;
#400 value1=32'd3608;value2=32'd3622;
#400 value1=32'd3638;value2=32'd3652;
#400 value1=32'd3668;value2=32'd3682;
#400 value1=32'd3698;value2=32'd3712;
#400 value1=32'd3728;value2=32'd3742;
#400 value1=32'd3758;value2=32'd3772;
#400 value1=32'd3788;value2=32'd3804;
#400 value1=32'd3818;value2=32'd3834;
#400 value1=32'd3848;value2=32'd3862;
#400 value1=32'd3874;value2=32'd3890;
#400 value1=32'd3904;value2=32'd3918;
#400 value1=32'd3934;value2=32'd3950;
#400 value1=32'd3966;value2=32'd3982;
#400 value1=32'd3998;value2=32'd4014;
#400 value1=32'd4032;value2=32'd4050;
#400 value1=32'd4064;value2=32'd4080;
#400 value1=32'd4096;value2=32'd4110;
#400 value1=32'd4124;value2=32'd4142;
#400 value1=32'd4160;value2=32'd4176;
#400 value1=32'd4192;value2=32'd4208;
#400 value1=32'd4224;value2=32'd4242;
#400 value1=32'd4260;value2=32'd4276;
#400 value1=32'd4292;value2=32'd4308;
#400 value1=32'd4322;value2=32'd4338;
#400 value1=32'd4356;value2=32'd4372;
#400 value1=32'd4390;value2=32'd4406;
#400 value1=32'd4422;value2=32'd4440;
#400 value1=32'd4456;value2=32'd4474;
#400 value1=32'd4490;value2=32'd4504;
#400 value1=32'd4522;value2=32'd4538;
#400 value1=32'd4556;value2=32'd4572;
#400 value1=32'd4590;value2=32'd4606;
#400 value1=32'd4624;value2=32'd4640;
#400 value1=32'd4652;value2=32'd4668;
#400 value1=32'd4682;value2=32'd4698;
#400 value1=32'd4712;value2=32'd4726;
#400 value1=32'd4742;value2=32'd4756;
#400 value1=32'd4772;value2=32'd4788;
#400 value1=32'd4802;value2=32'd4818;
#400 value1=32'd4832;value2=32'd4848;
#400 value1=32'd4862;value2=32'd4878;
#400 value1=32'd4892;value2=32'd4906;
#400 value1=32'd4922;value2=32'd4938;
#400 value1=32'd4954;value2=32'd4970;
#400 value1=32'd4988;value2=32'd5006;
#400 value1=32'd5022;value2=32'd5034;
#400 value1=32'd5048;value2=32'd5062;
#400 value1=32'd5078;value2=32'd5094;
#400 value1=32'd5108;value2=32'd5126;
#400 value1=32'd5144;value2=32'd5160;
#400 value1=32'd5176;value2=32'd5192;
#400 value1=32'd5208;value2=32'd5222;
#400 value1=32'd5236;value2=32'd5252;
#400 value1=32'd5268;value2=32'd5286;
#400 value1=32'd5304;value2=32'd5320;
#400 value1=32'd5336;value2=32'd5350;
#400 value1=32'd5364;value2=32'd5380;
#400 value1=32'd5396;value2=32'd5412;
#400 value1=32'd5428;value2=32'd5442;
#400 value1=32'd5456;value2=32'd5470;
#400 value1=32'd5484;value2=32'd5498;
#400 value1=32'd5514;value2=32'd5530;
#400 value1=32'd5546;value2=32'd5562;
#400 value1=32'd5574;value2=32'd5590;
#400 value1=32'd5602;value2=32'd5618;
#400 value1=32'd5636;value2=32'd5654;
#400 value1=32'd5672;value2=32'd5690;
#400 value1=32'd5706;value2=32'd5722;
#400 value1=32'd5738;value2=32'd5754;
#400 value1=32'd5770;value2=32'd5786;
#400 value1=32'd5804;value2=32'd5818;
#400 value1=32'd5834;value2=32'd5850;
#400 value1=32'd5868;value2=32'd5886;
#400 value1=32'd5902;value2=32'd5916;
#400 value1=32'd5932;value2=32'd5948;
#400 value1=32'd5966;value2=32'd5982;
#400 value1=32'd5998;value2=32'd6016;
#400 value1=32'd6030;value2=32'd6046;
#400 value1=32'd6062;value2=32'd6080;
#400 value1=32'd6094;value2=32'd6110;
#400 value1=32'd6124;value2=32'd6136;
#400 value1=32'd6152;value2=32'd6168;
#400 value1=32'd6184;value2=32'd6198;
#400 value1=32'd6212;value2=32'd6230;
#400 value1=32'd6248;value2=32'd6266;
#400 value1=32'd6284;value2=32'd6300;
#400 value1=32'd6316;value2=32'd6332;
#400 value1=32'd6348;value2=32'd6364;
#400 value1=32'd6380;value2=32'd6396;
#400 value1=32'd6412;value2=32'd6428;
#400 value1=32'd6440;value2=32'd6456;
#400 value1=32'd6468;value2=32'd6484;
#400 value1=32'd6500;value2=32'd6518;
#400 value1=32'd6534;value2=32'd6548;
#400 value1=32'd6566;value2=32'd6582;
#400 value1=32'd6600;value2=32'd6616;
#400 value1=32'd6632;value2=32'd6646;
#400 value1=32'd6664;value2=32'd6680;
#400 value1=32'd6696;value2=32'd6714;
#400 value1=32'd6730;value2=32'd6746;
#400 value1=32'd6760;value2=32'd6778;
#400 value1=32'd6794;value2=32'd6810;
#400 value1=32'd6824;value2=32'd6838;
#400 value1=32'd6854;value2=32'd6870;
#400 value1=32'd6886;value2=32'd6898;
#400 value1=32'd6912;value2=32'd6928;
#400 value1=32'd6944;value2=32'd6960;
#400 value1=32'd6976;value2=32'd6990;
#400 value1=32'd7004;value2=32'd7018;
#400 value1=32'd7032;value2=32'd7048;
#400 value1=32'd7064;value2=32'd7082;
#400 value1=32'd7096;value2=32'd7112;
#400 value1=32'd7128;value2=32'd7146;
#400 value1=32'd7164;value2=32'd7180;
#400 value1=32'd7194;value2=32'd7210;
#400 value1=32'd7226;value2=32'd7244;
#400 value1=32'd7260;value2=32'd7276;
#400 value1=32'd7294;value2=32'd7308;
#400 value1=32'd7324;value2=32'd7340;
#400 value1=32'd7358;value2=32'd7372;
#400 value1=32'd7388;value2=32'd7402;
#400 value1=32'd7414;value2=32'd7430;
#400 value1=32'd7446;value2=32'd7462;
#400 value1=32'd7476;value2=32'd7492;
#400 value1=32'd7508;value2=32'd7526;
#400 value1=32'd7542;value2=32'd7556;
#400 value1=32'd7574;value2=32'd7590;
#400 value1=32'd7608;value2=32'd7624;
#400 value1=32'd7640;value2=32'd7654;
#400 value1=32'd7672;value2=32'd7688;
#400 value1=32'd7704;value2=32'd7722;
#400 value1=32'd7738;value2=32'd7754;
#400 value1=32'd7768;value2=32'd7786;
#400 value1=32'd7802;value2=32'd7818;
#400 value1=32'd7832;value2=32'd7846;
#400 value1=32'd7862;value2=32'd7878;
#400 value1=32'd7894;value2=32'd7906;
#400 value1=32'd7920;value2=32'd7934;
#400 value1=32'd7948;value2=32'd7960;
#400 value1=32'd7972;value2=32'd7988;
#400 value1=32'd8004;value2=32'd8018;
#400 value1=32'd8032;value2=32'd8046;
#400 value1=32'd8060;value2=32'd8074;
#400 value1=32'd8090;value2=32'd8106;
#400 value1=32'd8122;value2=32'd8138;
#400 value1=32'd8150;value2=32'd8164;
#400 value1=32'd8180;value2=32'd8196;
#400 value1=32'd8210;value2=32'd8226;
#400 value1=32'd8240;value2=32'd8256;
#400 value1=32'd8272;value2=32'd8288;
#400 value1=32'd8304;value2=32'd8318;
#400 value1=32'd8332;value2=32'd8346;
#400 value1=32'd8360;value2=32'd8372;
#400 value1=32'd8386;value2=32'd8402;
#400 value1=32'd8418;value2=32'd8432;
#400 value1=32'd8448;value2=32'd8464;
#400 value1=32'd8480;value2=32'd8492;
#400 value1=32'd8504;value2=32'd8520;
#400 value1=32'd8534;value2=32'd8550;
#400 value1=32'd8566;value2=32'd8580;
#400 value1=32'd8592;value2=32'd8608;
#400 value1=32'd8622;value2=32'd8638;
#400 value1=32'd8654;value2=32'd8668;
#400 value1=32'd8680;value2=32'd8694;
#400 value1=32'd8708;value2=32'd8722;
#400 value1=32'd8736;value2=32'd0;
// dense
#400 value1=1;value2=1;
/*
*/

end

initial begin
#3608184 value1=0;value2=1;
#400 value1=2;value2=3;
#400 value1=4;value2=5;
#400 value1=6;value2=7;
#400 value1=8;value2=9;
#400 value1=10;value2=11;
#400 value1=12;value2=13;
#400 value1=14;value2=15;
#400 value1=16;value2=17;
#400 value1=18;value2=19;
#400 value1=20;value2=21;
#400 value1=22;value2=23;
#400 value1=24;value2=25;
#400 value1=26;value2=27;
#400 value1=28;value2=29;
#400 value1=30;value2=31;
#400 value1=32;value2=33;
#400 value1=34;value2=35;
#400 value1=36;value2=37;
#400 value1=38;value2=39;
#400 value1=40;value2=41;
#400 value1=42;value2=43;
#400 value1=44;value2=45;
#400 value1=46;value2=47;
#400 value1=48;value2=49;
#400 value1=50;value2=51;
#400 value1=52;value2=53;
#400 value1=54;value2=55;
#400 value1=56;value2=57;
#400 value1=58;value2=59;
#400 value1=60;value2=61;
#400 value1=62;value2=63;
#400 value1=64;value2=65;
#400 value1=66;value2=67;
#400 value1=68;value2=69;
#400 value1=70;value2=71;
#400 value1=72;value2=73;
#400 value1=74;value2=75;
#400 value1=76;value2=77;
#400 value1=78;value2=79;
#400 value1=80;value2=81;
#400 value1=82;value2=83;
#400 value1=84;value2=85;
#400 value1=86;value2=87;
#400 value1=88;value2=89;
#400 value1=90;value2=91;
#400 value1=92;value2=93;
#400 value1=94;value2=95;
#400 value1=96;value2=97;
#400 value1=98;value2=99;
#400 value1=100;value2=101;
#400 value1=102;value2=103;
#400 value1=104;value2=105;
#400 value1=106;value2=107;
#400 value1=108;value2=109;
#400 value1=110;value2=111;
#400 value1=112;value2=113;
#400 value1=114;value2=115;
#400 value1=116;value2=117;
#400 value1=118;value2=119;
#400 value1=120;value2=121;
#400 value1=122;value2=123;
#400 value1=124;value2=125;
#400 value1=126;value2=127;
#400 value1=128;value2=129;
#400 value1=130;value2=131;
#400 value1=132;value2=133;
#400 value1=134;value2=135;
#400 value1=136;value2=137;
#400 value1=138;value2=139;
#400 value1=140;value2=141;
#400 value1=142;value2=143;
#400 value1=144;value2=145;
#400 value1=146;value2=147;
#400 value1=148;value2=149;
#400 value1=150;value2=151;
#400 value1=152;value2=153;
#400 value1=154;value2=155;
#400 value1=156;value2=157;
#400 value1=158;value2=159;
#400 value1=160;value2=161;
#400 value1=162;value2=163;
#400 value1=164;value2=165;
#400 value1=166;value2=167;
#400 value1=168;value2=169;
#400 value1=170;value2=171;
#400 value1=172;value2=173;
#400 value1=174;value2=175;
#400 value1=176;value2=177;
#400 value1=178;value2=179;
#400 value1=180;value2=181;
#400 value1=182;value2=183;
#400 value1=184;value2=185;
#400 value1=186;value2=187;
#400 value1=188;value2=189;
#400 value1=190;value2=191;
#400 value1=192;value2=193;
#400 value1=194;value2=195;
#400 value1=196;value2=197;
#400 value1=198;value2=199;
#400 value1=200;value2=201;
#400 value1=202;value2=203;
#400 value1=204;value2=205;
#400 value1=206;value2=207;
#400 value1=208;value2=209;
#400 value1=210;value2=211;
#400 value1=212;value2=213;
#400 value1=214;value2=215;
#400 value1=216;value2=217;
#400 value1=218;value2=219;
#400 value1=220;value2=221;
#400 value1=222;value2=223;
#400 value1=224;value2=225;
#400 value1=226;value2=227;
#400 value1=228;value2=229;
#400 value1=230;value2=231;
#400 value1=232;value2=233;
#400 value1=234;value2=235;
#400 value1=236;value2=237;
#400 value1=238;value2=239;
#400 value1=240;value2=241;
#400 value1=242;value2=243;
#400 value1=244;value2=245;
#400 value1=246;value2=247;
#400 value1=248;value2=249;
#400 value1=250;value2=251;
#400 value1=252;value2=253;
#400 value1=254;value2=255;
#400 value1=256;value2=257;
#400 value1=258;value2=259;
#400 value1=260;value2=261;
#400 value1=262;value2=263;
#400 value1=264;value2=265;
#400 value1=266;value2=267;
#400 value1=268;value2=269;
#400 value1=270;value2=271;
#400 value1=272;value2=273;
#400 value1=274;value2=275;
#400 value1=276;value2=277;
#400 value1=278;value2=279;
#400 value1=280;value2=281;
#400 value1=282;value2=283;
#400 value1=284;value2=285;
#400 value1=286;value2=287;
#400 value1=288;value2=289;
#400 value1=290;value2=291;
#400 value1=292;value2=293;
#400 value1=294;value2=295;
#400 value1=296;value2=297;
#400 value1=298;value2=299;
#400 value1=300;value2=301;
#400 value1=302;value2=303;
#400 value1=304;value2=305;
#400 value1=306;value2=307;
#400 value1=308;value2=309;
#400 value1=310;value2=311;
#400 value1=312;value2=313;
#400 value1=314;value2=315;
#400 value1=316;value2=317;
#400 value1=318;value2=319;
#400 value1=320;value2=321;
#400 value1=322;value2=323;
#400 value1=324;value2=325;
#400 value1=326;value2=327;
#400 value1=328;value2=329;
#400 value1=330;value2=331;
#400 value1=332;value2=333;
#400 value1=334;value2=335;
#400 value1=336;value2=337;
#400 value1=338;value2=339;
#400 value1=340;value2=341;
#400 value1=342;value2=343;
#400 value1=344;value2=345;
#400 value1=346;value2=347;
#400 value1=348;value2=349;
#400 value1=350;value2=351;
#400 value1=352;value2=353;
#400 value1=354;value2=355;
#400 value1=356;value2=357;
#400 value1=358;value2=359;
#400 value1=360;value2=361;
#400 value1=362;value2=363;
#400 value1=364;value2=365;
#400 value1=366;value2=367;
#400 value1=368;value2=369;
#400 value1=370;value2=371;
#400 value1=372;value2=373;
#400 value1=374;value2=375;
#400 value1=376;value2=377;
#400 value1=378;value2=379;
#400 value1=380;value2=381;
#400 value1=382;value2=383;
#400 value1=384;value2=385;
#400 value1=386;value2=387;
#400 value1=388;value2=389;
#400 value1=390;value2=391;
#400 value1=392;value2=393;
#400 value1=394;value2=395;
#400 value1=396;value2=397;
#400 value1=398;value2=399;
#400 value1=400;value2=401;
#400 value1=402;value2=403;
#400 value1=404;value2=405;
#400 value1=406;value2=407;
#400 value1=408;value2=409;
#400 value1=410;value2=411;
#400 value1=412;value2=413;
#400 value1=414;value2=415;
#400 value1=416;value2=417;
#400 value1=418;value2=419;
#400 value1=420;value2=421;
#400 value1=422;value2=423;
#400 value1=424;value2=425;
#400 value1=426;value2=427;
#400 value1=428;value2=429;
#400 value1=430;value2=431;
#400 value1=432;value2=433;
#400 value1=434;value2=435;
#400 value1=436;value2=437;
#400 value1=438;value2=439;
#400 value1=440;value2=441;
#400 value1=442;value2=443;
#400 value1=444;value2=445;
#400 value1=446;value2=447;
#400 value1=448;value2=449;
#400 value1=450;value2=451;
#400 value1=452;value2=453;
#400 value1=454;value2=455;
#400 value1=456;value2=457;
#400 value1=458;value2=459;
#400 value1=460;value2=461;
#400 value1=462;value2=463;
#400 value1=464;value2=465;
#400 value1=466;value2=467;
#400 value1=468;value2=469;
#400 value1=470;value2=471;
#400 value1=472;value2=473;
#400 value1=474;value2=475;
#400 value1=476;value2=477;
#400 value1=478;value2=479;
#400 value1=480;value2=481;
#400 value1=482;value2=483;
#400 value1=484;value2=485;
#400 value1=486;value2=487;
#400 value1=488;value2=489;
#400 value1=490;value2=491;
#400 value1=492;value2=493;
#400 value1=494;value2=495;
#400 value1=496;value2=497;
#400 value1=498;value2=499;
#400 value1=500;value2=501;
#400 value1=502;value2=503;
#400 value1=504;value2=505;
#400 value1=506;value2=507;
#400 value1=508;value2=509;
#400 value1=510;value2=511;
#400 value1=512;value2=513;
#400 value1=514;value2=515;
#400 value1=516;value2=517;
#400 value1=518;value2=519;
#400 value1=520;value2=521;
#400 value1=522;value2=523;
#400 value1=524;value2=525;
#400 value1=526;value2=527;
#400 value1=528;value2=529;
#400 value1=530;value2=531;
#400 value1=532;value2=533;
#400 value1=534;value2=535;
#400 value1=536;value2=537;
#400 value1=538;value2=539;
#400 value1=540;value2=541;
#400 value1=542;value2=543;
#400 value1=544;value2=545;
#400 value1=546;value2=547;
#400 value1=548;value2=549;
#400 value1=550;value2=551;
#400 value1=552;value2=553;
#400 value1=554;value2=555;
#400 value1=556;value2=557;
#400 value1=558;value2=559;

#34 value1=0;value2=1;
#400 value1=2;value2=3;
#400 value1=4;value2=5;
#400 value1=6;value2=7;
#400 value1=8;value2=9;
#400 value1=10;value2=11;
#400 value1=12;value2=13;
#400 value1=14;value2=15;
#400 value1=16;value2=17;
#400 value1=18;value2=19;
#400 value1=20;value2=21;
#400 value1=22;value2=23;
#400 value1=24;value2=25;
#400 value1=26;value2=27;
#400 value1=28;value2=29;
#400 value1=30;value2=31;
#400 value1=32;value2=33;
#400 value1=34;value2=35;
#400 value1=36;value2=37;
#400 value1=38;value2=39;
#400 value1=40;value2=41;
#400 value1=42;value2=43;
#400 value1=44;value2=45;
#400 value1=46;value2=47;
#400 value1=48;value2=49;
#400 value1=50;value2=51;
#400 value1=52;value2=53;
#400 value1=54;value2=55;
#400 value1=56;value2=57;
#400 value1=58;value2=59;
#400 value1=60;value2=61;
#400 value1=62;value2=63;
#400 value1=64;value2=65;
#400 value1=66;value2=67;
#400 value1=68;value2=69;
#400 value1=70;value2=71;
#400 value1=72;value2=73;
#400 value1=74;value2=75;
#400 value1=76;value2=77;
#400 value1=78;value2=79;
#400 value1=80;value2=81;
#400 value1=82;value2=83;
#400 value1=84;value2=85;
#400 value1=86;value2=87;
#400 value1=88;value2=89;
#400 value1=90;value2=91;
#400 value1=92;value2=93;
#400 value1=94;value2=95;
#400 value1=96;value2=97;
#400 value1=98;value2=99;
#400 value1=100;value2=101;
#400 value1=102;value2=103;
#400 value1=104;value2=105;
#400 value1=106;value2=107;
#400 value1=108;value2=109;
#400 value1=110;value2=111;
#400 value1=112;value2=113;
#400 value1=114;value2=115;
#400 value1=116;value2=117;
#400 value1=118;value2=119;
#400 value1=120;value2=121;
#400 value1=122;value2=123;
#400 value1=124;value2=125;
#400 value1=126;value2=127;
#400 value1=128;value2=129;
#400 value1=130;value2=131;
#400 value1=132;value2=133;
#400 value1=134;value2=135;
#400 value1=136;value2=137;
#400 value1=138;value2=139;
#400 value1=140;value2=141;
#400 value1=142;value2=143;
#400 value1=144;value2=145;
#400 value1=146;value2=147;
#400 value1=148;value2=149;
#400 value1=150;value2=151;
#400 value1=152;value2=153;
#400 value1=154;value2=155;
#400 value1=156;value2=157;
#400 value1=158;value2=159;
#400 value1=160;value2=161;
#400 value1=162;value2=163;
#400 value1=164;value2=165;
#400 value1=166;value2=167;
#400 value1=168;value2=169;
#400 value1=170;value2=171;
#400 value1=172;value2=173;
#400 value1=174;value2=175;
#400 value1=176;value2=177;
#400 value1=178;value2=179;
#400 value1=180;value2=181;
#400 value1=182;value2=183;
#400 value1=184;value2=185;
#400 value1=186;value2=187;
#400 value1=188;value2=189;
#400 value1=190;value2=191;
#400 value1=192;value2=193;
#400 value1=194;value2=195;
#400 value1=196;value2=197;
#400 value1=198;value2=199;
#400 value1=200;value2=201;
#400 value1=202;value2=203;
#400 value1=204;value2=205;
#400 value1=206;value2=207;
#400 value1=208;value2=209;
#400 value1=210;value2=211;
#400 value1=212;value2=213;
#400 value1=214;value2=215;
#400 value1=216;value2=217;
#400 value1=218;value2=219;
#400 value1=220;value2=221;
#400 value1=222;value2=223;
#400 value1=224;value2=225;
#400 value1=226;value2=227;
#400 value1=228;value2=229;
#400 value1=230;value2=231;
#400 value1=232;value2=233;
#400 value1=234;value2=235;
#400 value1=236;value2=237;
#400 value1=238;value2=239;
#400 value1=240;value2=241;
#400 value1=242;value2=243;
#400 value1=244;value2=245;
#400 value1=246;value2=247;
#400 value1=248;value2=249;
#400 value1=250;value2=251;
#400 value1=252;value2=253;
#400 value1=254;value2=255;
#400 value1=256;value2=257;
#400 value1=258;value2=259;
#400 value1=260;value2=261;
#400 value1=262;value2=263;
#400 value1=264;value2=265;
#400 value1=266;value2=267;
#400 value1=268;value2=269;
#400 value1=270;value2=271;
#400 value1=272;value2=273;
#400 value1=274;value2=275;
#400 value1=276;value2=277;
#400 value1=278;value2=279;
#400 value1=280;value2=281;
#400 value1=282;value2=283;
#400 value1=284;value2=285;
#400 value1=286;value2=287;
#400 value1=288;value2=289;
#400 value1=290;value2=291;
#400 value1=292;value2=293;
#400 value1=294;value2=295;
#400 value1=296;value2=297;
#400 value1=298;value2=299;
#400 value1=300;value2=301;
#400 value1=302;value2=303;
#400 value1=304;value2=305;
#400 value1=306;value2=307;
#400 value1=308;value2=309;
#400 value1=310;value2=311;
#400 value1=312;value2=313;
#400 value1=314;value2=315;
#400 value1=316;value2=317;
#400 value1=318;value2=319;
#400 value1=320;value2=321;
#400 value1=322;value2=323;
#400 value1=324;value2=325;
#400 value1=326;value2=327;
#400 value1=328;value2=329;
#400 value1=330;value2=331;
#400 value1=332;value2=333;
#400 value1=334;value2=335;
#400 value1=336;value2=337;
#400 value1=338;value2=339;
#400 value1=340;value2=341;
#400 value1=342;value2=343;
#400 value1=344;value2=345;
#400 value1=346;value2=347;
#400 value1=348;value2=349;
#400 value1=350;value2=351;
#400 value1=352;value2=353;
#400 value1=354;value2=355;
#400 value1=356;value2=357;
#400 value1=358;value2=359;
#400 value1=360;value2=361;
#400 value1=362;value2=363;
#400 value1=364;value2=365;
#400 value1=366;value2=367;
#400 value1=368;value2=369;
#400 value1=370;value2=371;
#400 value1=372;value2=373;
#400 value1=374;value2=375;
#400 value1=376;value2=377;
#400 value1=378;value2=379;
#400 value1=380;value2=381;
#400 value1=382;value2=383;
#400 value1=384;value2=385;
#400 value1=386;value2=387;
#400 value1=388;value2=389;
#400 value1=390;value2=391;
#400 value1=392;value2=393;
#400 value1=394;value2=395;
#400 value1=396;value2=397;
#400 value1=398;value2=399;
#400 value1=400;value2=401;
#400 value1=402;value2=403;
#400 value1=404;value2=405;
#400 value1=406;value2=407;
#400 value1=408;value2=409;
#400 value1=410;value2=411;
#400 value1=412;value2=413;
#400 value1=414;value2=415;
#400 value1=416;value2=417;
#400 value1=418;value2=419;
#400 value1=420;value2=421;
#400 value1=422;value2=423;
#400 value1=424;value2=425;
#400 value1=426;value2=427;
#400 value1=428;value2=429;
#400 value1=430;value2=431;
#400 value1=432;value2=433;
#400 value1=434;value2=435;
#400 value1=436;value2=437;
#400 value1=438;value2=439;
#400 value1=440;value2=441;
#400 value1=442;value2=443;
#400 value1=444;value2=445;
#400 value1=446;value2=447;
#400 value1=448;value2=449;
#400 value1=450;value2=451;
#400 value1=452;value2=453;
#400 value1=454;value2=455;
#400 value1=456;value2=457;
#400 value1=458;value2=459;
#400 value1=460;value2=461;
#400 value1=462;value2=463;
#400 value1=464;value2=465;
#400 value1=466;value2=467;
#400 value1=468;value2=469;
#400 value1=470;value2=471;
#400 value1=472;value2=473;
#400 value1=474;value2=475;
#400 value1=476;value2=477;
#400 value1=478;value2=479;
#400 value1=480;value2=481;
#400 value1=482;value2=483;
#400 value1=484;value2=485;
#400 value1=486;value2=487;
#400 value1=488;value2=489;
#400 value1=490;value2=491;
#400 value1=492;value2=493;
#400 value1=494;value2=495;
#400 value1=496;value2=497;
#400 value1=498;value2=499;
#400 value1=500;value2=501;
#400 value1=502;value2=503;
#400 value1=504;value2=505;
#400 value1=506;value2=507;
#400 value1=508;value2=509;
#400 value1=510;value2=511;
#400 value1=512;value2=513;
#400 value1=514;value2=515;
#400 value1=516;value2=517;
#400 value1=518;value2=519;
#400 value1=520;value2=521;
#400 value1=522;value2=523;
#400 value1=524;value2=525;
#400 value1=526;value2=527;
#400 value1=528;value2=529;
#400 value1=530;value2=531;
#400 value1=532;value2=533;
#400 value1=534;value2=535;
#400 value1=536;value2=537;
#400 value1=538;value2=539;
#400 value1=540;value2=541;
#400 value1=542;value2=543;
#400 value1=544;value2=545;
#400 value1=546;value2=547;
#400 value1=548;value2=549;
#400 value1=550;value2=551;
#400 value1=552;value2=553;
#400 value1=554;value2=555;
#400 value1=556;value2=557;
#400 value1=558;value2=559;
end

initial begin
//value
#982154270 value1=32'd1;value2=32'd1;
#1747200 value1=32'd1;value2=32'd1;
//column
#400 value1=32'd1;value2=32'd4;
#400 value1=32'd5;value2=32'd6;
#400 value1=32'd8;value2=32'd14;
#400 value1=32'd15;value2=32'd16;
#400 value1=32'd20;value2=32'd22;
#400 value1=32'd106;value2=32'd107;
#400 value1=32'd110;value2=32'd112;
#400 value1=32'd0;value2=32'd4;
#400 value1=32'd5;value2=32'd7;
#400 value1=32'd9;value2=32'd27;
#400 value1=32'd28;value2=32'd32;
#400 value1=32'd34;value2=32'd105;
#400 value1=32'd118;value2=32'd119;
#400 value1=32'd122;value2=32'd124;
#400 value1=32'd3;value2=32'd4;
#400 value1=32'd10;value2=32'd12;
#400 value1=32'd27;value2=32'd39;
#400 value1=32'd43;value2=32'd45;
#400 value1=32'd106;value2=32'd130;
#400 value1=32'd133;value2=32'd135;
#400 value1=32'd2;value2=32'd5;
#400 value1=32'd11;value2=32'd13;
#400 value1=32'd28;value2=32'd39;
#400 value1=32'd53;value2=32'd55;
#400 value1=32'd107;value2=32'd130;
#400 value1=32'd143;value2=32'd145;
#400 value1=32'd0;value2=32'd1;
#400 value1=32'd2;value2=32'd5;
#400 value1=32'd10;value2=32'd12;
#400 value1=32'd29;value2=32'd40;
#400 value1=32'd50;value2=32'd62;
#400 value1=32'd64;value2=32'd108;
#400 value1=32'd131;value2=32'd141;
#400 value1=32'd152;value2=32'd154;
#400 value1=32'd0;value2=32'd1;
#400 value1=32'd3;value2=32'd4;
#400 value1=32'd11;value2=32'd13;
#400 value1=32'd30;value2=32'd41;
#400 value1=32'd51;value2=32'd70;
#400 value1=32'd72;value2=32'd109;
#400 value1=32'd132;value2=32'd142;
#400 value1=32'd160;value2=32'd162;
#400 value1=32'd0;value2=32'd7;
#400 value1=32'd8;value2=32'd10;
#400 value1=32'd11;value2=32'd31;
#400 value1=32'd42;value2=32'd52;
#400 value1=32'd77;value2=32'd79;
#400 value1=32'd110;value2=32'd133;
#400 value1=32'd143;value2=32'd169;
#400 value1=32'd1;value2=32'd6;
#400 value1=32'd9;value2=32'd10;
#400 value1=32'd11;value2=32'd32;
#400 value1=32'd43;value2=32'd53;
#400 value1=32'd85;value2=32'd111;
#400 value1=32'd134;value2=32'd144;
#400 value1=32'd168;value2=32'd175;
#400 value1=32'd0;value2=32'd6;
#400 value1=32'd9;value2=32'd12;
#400 value1=32'd13;value2=32'd33;
#400 value1=32'd44;value2=32'd54;
#400 value1=32'd84;value2=32'd90;
#400 value1=32'd112;value2=32'd135;
#400 value1=32'd145;value2=32'd169;
#400 value1=32'd1;value2=32'd7;
#400 value1=32'd8;value2=32'd12;
#400 value1=32'd13;value2=32'd34;
#400 value1=32'd45;value2=32'd55;
#400 value1=32'd85;value2=32'd113;
#400 value1=32'd136;value2=32'd146;
#400 value1=32'd170;value2=32'd181;
#400 value1=32'd2;value2=32'd4;
#400 value1=32'd6;value2=32'd7;
#400 value1=32'd11;value2=32'd12;
#400 value1=32'd35;value2=32'd46;
#400 value1=32'd56;value2=32'd86;
#400 value1=32'd95;value2=32'd114;
#400 value1=32'd137;value2=32'd147;
#400 value1=32'd171;value2=32'd182;
#400 value1=32'd3;value2=32'd5;
#400 value1=32'd6;value2=32'd7;
#400 value1=32'd10;value2=32'd13;
#400 value1=32'd36;value2=32'd47;
#400 value1=32'd57;value2=32'd87;
#400 value1=32'd96;value2=32'd115;
#400 value1=32'd138;value2=32'd148;
#400 value1=32'd172;value2=32'd183;
#400 value1=32'd2;value2=32'd4;
#400 value1=32'd8;value2=32'd9;
#400 value1=32'd10;value2=32'd13;
#400 value1=32'd37;value2=32'd48;
#400 value1=32'd58;value2=32'd88;
#400 value1=32'd97;value2=32'd116;
#400 value1=32'd139;value2=32'd149;
#400 value1=32'd173;value2=32'd184;
#400 value1=32'd3;value2=32'd5;
#400 value1=32'd8;value2=32'd9;
#400 value1=32'd11;value2=32'd12;
#400 value1=32'd38;value2=32'd49;
#400 value1=32'd59;value2=32'd89;
#400 value1=32'd98;value2=32'd117;
#400 value1=32'd140;value2=32'd150;
#400 value1=32'd174;value2=32'd185;
#400 value1=32'd0;value2=32'd17;
#400 value1=32'd18;value2=32'd20;
#400 value1=32'd22;value2=32'd29;
#400 value1=32'd30;value2=32'd31;
#400 value1=32'd33;value2=32'd105;
#400 value1=32'd196;value2=32'd197;
#400 value1=32'd200;value2=32'd202;
#400 value1=32'd0;value2=32'd16;
#400 value1=32'd17;value2=32'd23;
#400 value1=32'd25;value2=32'd27;
#400 value1=32'd40;value2=32'd41;
#400 value1=32'd42;value2=32'd44;
#400 value1=32'd106;value2=32'd208;
#400 value1=32'd211;value2=32'd213;
#400 value1=32'd0;value2=32'd15;
#400 value1=32'd18;value2=32'd24;
#400 value1=32'd26;value2=32'd28;
#400 value1=32'd50;value2=32'd51;
#400 value1=32'd52;value2=32'd54;
#400 value1=32'd107;value2=32'd208;
#400 value1=32'd221;value2=32'd223;
#400 value1=32'd14;value2=32'd15;
#400 value1=32'd18;value2=32'd23;
#400 value1=32'd25;value2=32'd29;
#400 value1=32'd60;value2=32'd61;
#400 value1=32'd63;value2=32'd108;
#400 value1=32'd209;value2=32'd219;
#400 value1=32'd230;value2=32'd232;
#400 value1=32'd14;value2=32'd16;
#400 value1=32'd17;value2=32'd24;
#400 value1=32'd26;value2=32'd30;
#400 value1=32'd60;value2=32'd69;
#400 value1=32'd71;value2=32'd109;
#400 value1=32'd210;value2=32'd220;
#400 value1=32'd238;value2=32'd240;
#400 value1=32'd20;value2=32'd21;
#400 value1=32'd23;value2=32'd24;
#400 value1=32'd31;value2=32'd61;
#400 value1=32'd69;value2=32'd78;
#400 value1=32'd110;value2=32'd211;
#400 value1=32'd221;value2=32'd247;
#400 value1=32'd0;value2=32'd14;
#400 value1=32'd19;value2=32'd22;
#400 value1=32'd23;value2=32'd24;
#400 value1=32'd32;value2=32'd62;
#400 value1=32'd70;value2=32'd77;
#400 value1=32'd84;value2=32'd111;
#400 value1=32'd212;value2=32'd222;
#400 value1=32'd246;value2=32'd253;
#400 value1=32'd19;value2=32'd22;
#400 value1=32'd25;value2=32'd26;
#400 value1=32'd33;value2=32'd63;
#400 value1=32'd71;value2=32'd78;
#400 value1=32'd112;value2=32'd213;
#400 value1=32'd223;value2=32'd247;
#400 value1=32'd0;value2=32'd14;
#400 value1=32'd20;value2=32'd21;
#400 value1=32'd25;value2=32'd26;
#400 value1=32'd34;value2=32'd64;
#400 value1=32'd72;value2=32'd79;
#400 value1=32'd90;value2=32'd113;
#400 value1=32'd214;value2=32'd224;
#400 value1=32'd248;value2=32'd259;
#400 value1=32'd15;value2=32'd17;
#400 value1=32'd19;value2=32'd20;
#400 value1=32'd24;value2=32'd25;
#400 value1=32'd35;value2=32'd65;
#400 value1=32'd73;value2=32'd80;
#400 value1=32'd91;value2=32'd114;
#400 value1=32'd215;value2=32'd225;
#400 value1=32'd249;value2=32'd260;
#400 value1=32'd16;value2=32'd18;
#400 value1=32'd19;value2=32'd20;
#400 value1=32'd23;value2=32'd26;
#400 value1=32'd36;value2=32'd66;
#400 value1=32'd74;value2=32'd81;
#400 value1=32'd92;value2=32'd115;
#400 value1=32'd216;value2=32'd226;
#400 value1=32'd250;value2=32'd261;
#400 value1=32'd15;value2=32'd17;
#400 value1=32'd21;value2=32'd22;
#400 value1=32'd23;value2=32'd26;
#400 value1=32'd37;value2=32'd67;
#400 value1=32'd75;value2=32'd82;
#400 value1=32'd93;value2=32'd116;
#400 value1=32'd217;value2=32'd227;
#400 value1=32'd251;value2=32'd262;
#400 value1=32'd16;value2=32'd18;
#400 value1=32'd21;value2=32'd22;
#400 value1=32'd24;value2=32'd25;
#400 value1=32'd38;value2=32'd68;
#400 value1=32'd76;value2=32'd83;
#400 value1=32'd94;value2=32'd117;
#400 value1=32'd218;value2=32'd228;
#400 value1=32'd252;value2=32'd263;
#400 value1=32'd1;value2=32'd2;
#400 value1=32'd15;value2=32'd28;
#400 value1=32'd29;value2=32'd35;
#400 value1=32'd37;value2=32'd40;
#400 value1=32'd41;value2=32'd43;
#400 value1=32'd45;value2=32'd118;
#400 value1=32'd196;value2=32'd274;
#400 value1=32'd277;value2=32'd279;
#400 value1=32'd1;value2=32'd3;
#400 value1=32'd16;value2=32'd27;
#400 value1=32'd30;value2=32'd36;
#400 value1=32'd38;value2=32'd50;
#400 value1=32'd51;value2=32'd53;
#400 value1=32'd55;value2=32'd119;
#400 value1=32'd197;value2=32'd274;
#400 value1=32'd287;value2=32'd289;
#400 value1=32'd4;value2=32'd14;
#400 value1=32'd17;value2=32'd27;
#400 value1=32'd30;value2=32'd35;
#400 value1=32'd37;value2=32'd60;
#400 value1=32'd62;value2=32'd64;
#400 value1=32'd120;value2=32'd198;
#400 value1=32'd275;value2=32'd285;
#400 value1=32'd296;value2=32'd298;
#400 value1=32'd5;value2=32'd14;
#400 value1=32'd18;value2=32'd28;
#400 value1=32'd29;value2=32'd36;
#400 value1=32'd38;value2=32'd60;
#400 value1=32'd70;value2=32'd72;
#400 value1=32'd121;value2=32'd199;
#400 value1=32'd276;value2=32'd286;
#400 value1=32'd304;value2=32'd306;
#400 value1=32'd6;value2=32'd14;
#400 value1=32'd19;value2=32'd32;
#400 value1=32'd33;value2=32'd35;
#400 value1=32'd36;value2=32'd61;
#400 value1=32'd69;value2=32'd77;
#400 value1=32'd79;value2=32'd122;
#400 value1=32'd200;value2=32'd277;
#400 value1=32'd287;value2=32'd313;
#400 value1=32'd1;value2=32'd7;
#400 value1=32'd20;value2=32'd31;
#400 value1=32'd34;value2=32'd35;
#400 value1=32'd36;value2=32'd62;
#400 value1=32'd70;value2=32'd85;
#400 value1=32'd123;value2=32'd201;
#400 value1=32'd278;value2=32'd288;
#400 value1=32'd312;value2=32'd319;
#400 value1=32'd8;value2=32'd14;
#400 value1=32'd21;value2=32'd31;
#400 value1=32'd34;value2=32'd37;
#400 value1=32'd38;value2=32'd63;
#400 value1=32'd71;value2=32'd84;
#400 value1=32'd90;value2=32'd124;
#400 value1=32'd202;value2=32'd279;
#400 value1=32'd289;value2=32'd313;
#400 value1=32'd1;value2=32'd9;
#400 value1=32'd22;value2=32'd32;
#400 value1=32'd33;value2=32'd37;
#400 value1=32'd38;value2=32'd64;
#400 value1=32'd72;value2=32'd85;
#400 value1=32'd125;value2=32'd203;
#400 value1=32'd280;value2=32'd290;
#400 value1=32'd314;value2=32'd325;
#400 value1=32'd10;value2=32'd23;
#400 value1=32'd27;value2=32'd29;
#400 value1=32'd31;value2=32'd32;
#400 value1=32'd36;value2=32'd37;
#400 value1=32'd65;value2=32'd73;
#400 value1=32'd86;value2=32'd95;
#400 value1=32'd126;value2=32'd204;
#400 value1=32'd281;value2=32'd291;
#400 value1=32'd315;value2=32'd326;
#400 value1=32'd11;value2=32'd24;
#400 value1=32'd28;value2=32'd30;
#400 value1=32'd31;value2=32'd32;
#400 value1=32'd35;value2=32'd38;
#400 value1=32'd66;value2=32'd74;
#400 value1=32'd87;value2=32'd96;
#400 value1=32'd127;value2=32'd205;
#400 value1=32'd282;value2=32'd292;
#400 value1=32'd316;value2=32'd327;
#400 value1=32'd12;value2=32'd25;
#400 value1=32'd27;value2=32'd29;
#400 value1=32'd33;value2=32'd34;
#400 value1=32'd35;value2=32'd38;
#400 value1=32'd67;value2=32'd75;
#400 value1=32'd88;value2=32'd97;
#400 value1=32'd128;value2=32'd206;
#400 value1=32'd283;value2=32'd293;
#400 value1=32'd317;value2=32'd328;
#400 value1=32'd13;value2=32'd26;
#400 value1=32'd28;value2=32'd30;
#400 value1=32'd33;value2=32'd34;
#400 value1=32'd36;value2=32'd37;
#400 value1=32'd68;value2=32'd76;
#400 value1=32'd89;value2=32'd98;
#400 value1=32'd129;value2=32'd207;
#400 value1=32'd284;value2=32'd294;
#400 value1=32'd318;value2=32'd329;
#400 value1=32'd2;value2=32'd3;
#400 value1=32'd41;value2=32'd47;
#400 value1=32'd49;value2=32'd50;
#400 value1=32'd56;value2=32'd58;
#400 value1=32'd130;value2=32'd208;
#400 value1=32'd342;value2=32'd344;
#400 value1=32'd4;value2=32'd15;
#400 value1=32'd27;value2=32'd41;
#400 value1=32'd46;value2=32'd48;
#400 value1=32'd50;value2=32'd65;
#400 value1=32'd67;value2=32'd131;
#400 value1=32'd209;value2=32'd340;
#400 value1=32'd351;value2=32'd353;
#400 value1=32'd5;value2=32'd15;
#400 value1=32'd27;value2=32'd39;
#400 value1=32'd40;value2=32'd47;
#400 value1=32'd49;value2=32'd51;
#400 value1=32'd60;value2=32'd73;
#400 value1=32'd75;value2=32'd132;
#400 value1=32'd210;value2=32'd341;
#400 value1=32'd359;value2=32'd361;
#400 value1=32'd6;value2=32'd15;
#400 value1=32'd43;value2=32'd44;
#400 value1=32'd46;value2=32'd47;
#400 value1=32'd52;value2=32'd61;
#400 value1=32'd80;value2=32'd82;
#400 value1=32'd133;value2=32'd211;
#400 value1=32'd342;value2=32'd368;
#400 value1=32'd2;value2=32'd7;
#400 value1=32'd27;value2=32'd42;
#400 value1=32'd45;value2=32'd46;
#400 value1=32'd47;value2=32'd53;
#400 value1=32'd62;value2=32'd86;
#400 value1=32'd88;value2=32'd134;
#400 value1=32'd212;value2=32'd343;
#400 value1=32'd367;value2=32'd374;
#400 value1=32'd8;value2=32'd15;
#400 value1=32'd42;value2=32'd45;
#400 value1=32'd48;value2=32'd49;
#400 value1=32'd54;value2=32'd63;
#400 value1=32'd91;value2=32'd93;
#400 value1=32'd135;value2=32'd213;
#400 value1=32'd344;value2=32'd368;
#400 value1=32'd2;value2=32'd9;
#400 value1=32'd27;value2=32'd43;
#400 value1=32'd44;value2=32'd48;
#400 value1=32'd49;value2=32'd55;
#400 value1=32'd64;value2=32'd95;
#400 value1=32'd97;value2=32'd136;
#400 value1=32'd214;value2=32'd345;
#400 value1=32'd369;value2=32'd380;
#400 value1=32'd10;value2=32'd40;
#400 value1=32'd42;value2=32'd43;
#400 value1=32'd47;value2=32'd48;
#400 value1=32'd56;value2=32'd65;
#400 value1=32'd100;value2=32'd137;
#400 value1=32'd215;value2=32'd346;
#400 value1=32'd370;value2=32'd381;
#400 value1=32'd11;value2=32'd39;
#400 value1=32'd41;value2=32'd42;
#400 value1=32'd43;value2=32'd46;
#400 value1=32'd49;value2=32'd57;
#400 value1=32'd66;value2=32'd99;
#400 value1=32'd102;value2=32'd138;
#400 value1=32'd216;value2=32'd347;
#400 value1=32'd371;value2=32'd382;
#400 value1=32'd12;value2=32'd40;
#400 value1=32'd44;value2=32'd45;
#400 value1=32'd46;value2=32'd49;
#400 value1=32'd58;value2=32'd67;
#400 value1=32'd100;value2=32'd139;
#400 value1=32'd217;value2=32'd348;
#400 value1=32'd372;value2=32'd383;
#400 value1=32'd13;value2=32'd39;
#400 value1=32'd41;value2=32'd44;
#400 value1=32'd45;value2=32'd47;
#400 value1=32'd48;value2=32'd59;
#400 value1=32'd68;value2=32'd101;
#400 value1=32'd104;value2=32'd140;
#400 value1=32'd218;value2=32'd349;
#400 value1=32'd373;value2=32'd384;
#400 value1=32'd4;value2=32'd16;
#400 value1=32'd28;value2=32'd39;
#400 value1=32'd40;value2=32'd51;
#400 value1=32'd56;value2=32'd58;
#400 value1=32'd60;value2=32'd66;
#400 value1=32'd68;value2=32'd141;
#400 value1=32'd219;value2=32'd340;
#400 value1=32'd396;value2=32'd398;
#400 value1=32'd5;value2=32'd16;
#400 value1=32'd28;value2=32'd41;
#400 value1=32'd50;value2=32'd57;
#400 value1=32'd59;value2=32'd74;
#400 value1=32'd76;value2=32'd142;
#400 value1=32'd220;value2=32'd341;
#400 value1=32'd404;value2=32'd406;
#400 value1=32'd6;value2=32'd16;
#400 value1=32'd42;value2=32'd53;
#400 value1=32'd54;value2=32'd56;
#400 value1=32'd57;value2=32'd69;
#400 value1=32'd81;value2=32'd83;
#400 value1=32'd143;value2=32'd221;
#400 value1=32'd342;value2=32'd413;
#400 value1=32'd3;value2=32'd7;
#400 value1=32'd28;value2=32'd43;
#400 value1=32'd52;value2=32'd55;
#400 value1=32'd56;value2=32'd57;
#400 value1=32'd70;value2=32'd87;
#400 value1=32'd89;value2=32'd144;
#400 value1=32'd222;value2=32'd343;
#400 value1=32'd412;value2=32'd419;
#400 value1=32'd8;value2=32'd16;
#400 value1=32'd44;value2=32'd52;
#400 value1=32'd55;value2=32'd58;
#400 value1=32'd59;value2=32'd71;
#400 value1=32'd92;value2=32'd94;
#400 value1=32'd145;value2=32'd223;
#400 value1=32'd344;value2=32'd413;
#400 value1=32'd3;value2=32'd9;
#400 value1=32'd28;value2=32'd45;
#400 value1=32'd53;value2=32'd54;
#400 value1=32'd58;value2=32'd59;
#400 value1=32'd72;value2=32'd96;
#400 value1=32'd98;value2=32'd146;
#400 value1=32'd224;value2=32'd345;
#400 value1=32'd414;value2=32'd425;
#400 value1=32'd10;value2=32'd39;
#400 value1=32'd46;value2=32'd50;
#400 value1=32'd52;value2=32'd53;
#400 value1=32'd57;value2=32'd58;
#400 value1=32'd73;value2=32'd99;
#400 value1=32'd101;value2=32'd147;
#400 value1=32'd225;value2=32'd346;
#400 value1=32'd415;value2=32'd426;
#400 value1=32'd11;value2=32'd47;
#400 value1=32'd51;value2=32'd52;
#400 value1=32'd53;value2=32'd56;
#400 value1=32'd59;value2=32'd74;
#400 value1=32'd103;value2=32'd148;
#400 value1=32'd226;value2=32'd347;
#400 value1=32'd416;value2=32'd427;
#400 value1=32'd12;value2=32'd39;
#400 value1=32'd48;value2=32'd50;
#400 value1=32'd54;value2=32'd55;
#400 value1=32'd56;value2=32'd59;
#400 value1=32'd75;value2=32'd102;
#400 value1=32'd104;value2=32'd149;
#400 value1=32'd227;value2=32'd348;
#400 value1=32'd417;value2=32'd428;
#400 value1=32'd13;value2=32'd49;
#400 value1=32'd51;value2=32'd54;
#400 value1=32'd55;value2=32'd57;
#400 value1=32'd58;value2=32'd76;
#400 value1=32'd103;value2=32'd150;
#400 value1=32'd228;value2=32'd349;
#400 value1=32'd418;value2=32'd429;
#400 value1=32'd17;value2=32'd18;
#400 value1=32'd29;value2=32'd30;
#400 value1=32'd41;value2=32'd50;
#400 value1=32'd66;value2=32'd68;
#400 value1=32'd73;value2=32'd75;
#400 value1=32'd151;value2=32'd229;
#400 value1=32'd350;value2=32'd395;
#400 value1=32'd440;value2=32'd442;
#400 value1=32'd17;value2=32'd19;
#400 value1=32'd31;value2=32'd42;
#400 value1=32'd62;value2=32'd63;
#400 value1=32'd65;value2=32'd66;
#400 value1=32'd69;value2=32'd80;
#400 value1=32'd82;value2=32'd152;
#400 value1=32'd230;value2=32'd351;
#400 value1=32'd396;value2=32'd449;
#400 value1=32'd4;value2=32'd20;
#400 value1=32'd29;value2=32'd32;
#400 value1=32'd43;value2=32'd61;
#400 value1=32'd64;value2=32'd65;
#400 value1=32'd66;value2=32'd70;
#400 value1=32'd86;value2=32'd88;
#400 value1=32'd153;value2=32'd231;
#400 value1=32'd352;value2=32'd397;
#400 value1=32'd448;value2=32'd455;
#400 value1=32'd17;value2=32'd21;
#400 value1=32'd33;value2=32'd44;
#400 value1=32'd61;value2=32'd64;
#400 value1=32'd67;value2=32'd68;
#400 value1=32'd71;value2=32'd91;
#400 value1=32'd93;value2=32'd154;
#400 value1=32'd232;value2=32'd353;
#400 value1=32'd398;value2=32'd449;
#400 value1=32'd4;value2=32'd22;
#400 value1=32'd29;value2=32'd34;
#400 value1=32'd45;value2=32'd62;
#400 value1=32'd63;value2=32'd67;
#400 value1=32'd68;value2=32'd72;
#400 value1=32'd95;value2=32'd97;
#400 value1=32'd155;value2=32'd233;
#400 value1=32'd354;value2=32'd399;
#400 value1=32'd450;value2=32'd461;
#400 value1=32'd23;value2=32'd35;
#400 value1=32'd40;value2=32'd46;
#400 value1=32'd61;value2=32'd62;
#400 value1=32'd66;value2=32'd67;
#400 value1=32'd73;value2=32'd100;
#400 value1=32'd156;value2=32'd234;
#400 value1=32'd355;value2=32'd400;
#400 value1=32'd451;value2=32'd462;
#400 value1=32'd24;value2=32'd36;
#400 value1=32'd47;value2=32'd50;
#400 value1=32'd60;value2=32'd61;
#400 value1=32'd62;value2=32'd65;
#400 value1=32'd68;value2=32'd74;
#400 value1=32'd99;value2=32'd102;
#400 value1=32'd157;value2=32'd235;
#400 value1=32'd356;value2=32'd401;
#400 value1=32'd452;value2=32'd463;
#400 value1=32'd25;value2=32'd37;
#400 value1=32'd40;value2=32'd48;
#400 value1=32'd63;value2=32'd64;
#400 value1=32'd65;value2=32'd68;
#400 value1=32'd75;value2=32'd100;
#400 value1=32'd158;value2=32'd236;
#400 value1=32'd357;value2=32'd402;
#400 value1=32'd453;value2=32'd464;
#400 value1=32'd26;value2=32'd38;
#400 value1=32'd49;value2=32'd50;
#400 value1=32'd60;value2=32'd63;
#400 value1=32'd64;value2=32'd66;
#400 value1=32'd67;value2=32'd76;
#400 value1=32'd101;value2=32'd104;
#400 value1=32'd159;value2=32'd237;
#400 value1=32'd358;value2=32'd403;
#400 value1=32'd454;value2=32'd465;
#400 value1=32'd18;value2=32'd19;
#400 value1=32'd31;value2=32'd52;
#400 value1=32'd61;value2=32'd70;
#400 value1=32'd71;value2=32'd73;
#400 value1=32'd74;value2=32'd81;
#400 value1=32'd83;value2=32'd160;
#400 value1=32'd238;value2=32'd359;
#400 value1=32'd404;value2=32'd477;
#400 value1=32'd5;value2=32'd20;
#400 value1=32'd30;value2=32'd32;
#400 value1=32'd53;value2=32'd62;
#400 value1=32'd69;value2=32'd72;
#400 value1=32'd73;value2=32'd74;
#400 value1=32'd87;value2=32'd89;
#400 value1=32'd161;value2=32'd239;
#400 value1=32'd360;value2=32'd405;
#400 value1=32'd476;value2=32'd483;
#400 value1=32'd18;value2=32'd21;
#400 value1=32'd33;value2=32'd54;
#400 value1=32'd63;value2=32'd69;
#400 value1=32'd72;value2=32'd75;
#400 value1=32'd76;value2=32'd92;
#400 value1=32'd94;value2=32'd162;
#400 value1=32'd240;value2=32'd361;
#400 value1=32'd406;value2=32'd477;
#400 value1=32'd5;value2=32'd22;
#400 value1=32'd30;value2=32'd34;
#400 value1=32'd55;value2=32'd64;
#400 value1=32'd70;value2=32'd71;
#400 value1=32'd75;value2=32'd76;
#400 value1=32'd96;value2=32'd98;
#400 value1=32'd163;value2=32'd241;
#400 value1=32'd362;value2=32'd407;
#400 value1=32'd478;value2=32'd489;
#400 value1=32'd23;value2=32'd35;
#400 value1=32'd41;value2=32'd56;
#400 value1=32'd60;value2=32'd65;
#400 value1=32'd69;value2=32'd70;
#400 value1=32'd74;value2=32'd75;
#400 value1=32'd99;value2=32'd101;
#400 value1=32'd164;value2=32'd242;
#400 value1=32'd363;value2=32'd408;
#400 value1=32'd479;value2=32'd490;
#400 value1=32'd24;value2=32'd36;
#400 value1=32'd51;value2=32'd57;
#400 value1=32'd66;value2=32'd69;
#400 value1=32'd70;value2=32'd73;
#400 value1=32'd76;value2=32'd103;
#400 value1=32'd165;value2=32'd243;
#400 value1=32'd364;value2=32'd409;
#400 value1=32'd480;value2=32'd491;
#400 value1=32'd25;value2=32'd37;
#400 value1=32'd41;value2=32'd58;
#400 value1=32'd60;value2=32'd67;
#400 value1=32'd71;value2=32'd72;
#400 value1=32'd73;value2=32'd76;
#400 value1=32'd102;value2=32'd104;
#400 value1=32'd166;value2=32'd244;
#400 value1=32'd365;value2=32'd410;
#400 value1=32'd481;value2=32'd492;
#400 value1=32'd26;value2=32'd38;
#400 value1=32'd51;value2=32'd59;
#400 value1=32'd68;value2=32'd71;
#400 value1=32'd72;value2=32'd74;
#400 value1=32'd75;value2=32'd103;
#400 value1=32'd167;value2=32'd245;
#400 value1=32'd366;value2=32'd411;
#400 value1=32'd482;value2=32'd493;
#400 value1=32'd6;value2=32'd20;
#400 value1=32'd31;value2=32'd79;
#400 value1=32'd80;value2=32'd81;
#400 value1=32'd84;value2=32'd86;
#400 value1=32'd87;value2=32'd168;
#400 value1=32'd246;value2=32'd367;
#400 value1=32'd412;value2=32'd504;
#400 value1=32'd19;value2=32'd21;
#400 value1=32'd79;value2=32'd82;
#400 value1=32'd83;value2=32'd84;
#400 value1=32'd91;value2=32'd92;
#400 value1=32'd169;value2=32'd247;
#400 value1=32'd368;value2=32'd413;
#400 value1=32'd6;value2=32'd22;
#400 value1=32'd31;value2=32'd77;
#400 value1=32'd78;value2=32'd82;
#400 value1=32'd83;value2=32'd85;
#400 value1=32'd90;value2=32'd95;
#400 value1=32'd96;value2=32'd170;
#400 value1=32'd248;value2=32'd369;
#400 value1=32'd414;value2=32'd510;
#400 value1=32'd23;value2=32'd42;
#400 value1=32'd61;value2=32'd77;
#400 value1=32'd81;value2=32'd82;
#400 value1=32'd86;value2=32'd91;
#400 value1=32'd99;value2=32'd171;
#400 value1=32'd249;value2=32'd370;
#400 value1=32'd415;value2=32'd511;
#400 value1=32'd24;value2=32'd52;
#400 value1=32'd69;value2=32'd77;
#400 value1=32'd80;value2=32'd83;
#400 value1=32'd87;value2=32'd92;
#400 value1=32'd99;value2=32'd172;
#400 value1=32'd250;value2=32'd371;
#400 value1=32'd416;value2=32'd512;
#400 value1=32'd25;value2=32'd42;
#400 value1=32'd61;value2=32'd78;
#400 value1=32'd79;value2=32'd80;
#400 value1=32'd83;value2=32'd88;
#400 value1=32'd93;value2=32'd100;
#400 value1=32'd102;value2=32'd173;
#400 value1=32'd251;value2=32'd372;
#400 value1=32'd417;value2=32'd513;
#400 value1=32'd26;value2=32'd52;
#400 value1=32'd69;value2=32'd78;
#400 value1=32'd79;value2=32'd81;
#400 value1=32'd82;value2=32'd89;
#400 value1=32'd94;value2=32'd101;
#400 value1=32'd103;value2=32'd174;
#400 value1=32'd252;value2=32'd373;
#400 value1=32'd418;value2=32'd514;
#400 value1=32'd8;value2=32'd20;
#400 value1=32'd33;value2=32'd77;
#400 value1=32'd78;value2=32'd85;
#400 value1=32'd88;value2=32'd89;
#400 value1=32'd90;value2=32'd91;
#400 value1=32'd92;value2=32'd175;
#400 value1=32'd253;value2=32'd374;
#400 value1=32'd419;value2=32'd504;
#400 value1=32'd7;value2=32'd9;
#400 value1=32'd32;value2=32'd34;
#400 value1=32'd79;value2=32'd84;
#400 value1=32'd88;value2=32'd89;
#400 value1=32'd95;value2=32'd96;
#400 value1=32'd176;value2=32'd254;
#400 value1=32'd375;value2=32'd420;
#400 value1=32'd505;value2=32'd525;
#400 value1=32'd10;value2=32'd35;
#400 value1=32'd43;value2=32'd62;
#400 value1=32'd77;value2=32'd80;
#400 value1=32'd87;value2=32'd88;
#400 value1=32'd95;value2=32'd99;
#400 value1=32'd177;value2=32'd255;
#400 value1=32'd376;value2=32'd421;
#400 value1=32'd506;value2=32'd526;
#400 value1=32'd11;value2=32'd36;
#400 value1=32'd53;value2=32'd70;
#400 value1=32'd77;value2=32'd81;
#400 value1=32'd86;value2=32'd89;
#400 value1=32'd96;value2=32'd99;
#400 value1=32'd178;value2=32'd256;
#400 value1=32'd377;value2=32'd422;
#400 value1=32'd507;value2=32'd527;
#400 value1=32'd12;value2=32'd37;
#400 value1=32'd43;value2=32'd62;
#400 value1=32'd82;value2=32'd84;
#400 value1=32'd85;value2=32'd86;
#400 value1=32'd89;value2=32'd97;
#400 value1=32'd100;value2=32'd102;
#400 value1=32'd179;value2=32'd257;
#400 value1=32'd378;value2=32'd423;
#400 value1=32'd508;value2=32'd528;
#400 value1=32'd13;value2=32'd38;
#400 value1=32'd53;value2=32'd70;
#400 value1=32'd83;value2=32'd84;
#400 value1=32'd85;value2=32'd87;
#400 value1=32'd88;value2=32'd98;
#400 value1=32'd101;value2=32'd103;
#400 value1=32'd180;value2=32'd258;
#400 value1=32'd379;value2=32'd424;
#400 value1=32'd509;value2=32'd529;
#400 value1=32'd8;value2=32'd22;
#400 value1=32'd33;value2=32'd79;
#400 value1=32'd84;value2=32'd93;
#400 value1=32'd94;value2=32'd97;
#400 value1=32'd98;value2=32'd181;
#400 value1=32'd259;value2=32'd380;
#400 value1=32'd425;value2=32'd510;
#400 value1=32'd23;value2=32'd44;
#400 value1=32'd63;value2=32'd78;
#400 value1=32'd80;value2=32'd84;
#400 value1=32'd92;value2=32'd93;
#400 value1=32'd95;value2=32'd100;
#400 value1=32'd101;value2=32'd182;
#400 value1=32'd260;value2=32'd381;
#400 value1=32'd426;value2=32'd511;
#400 value1=32'd24;value2=32'd54;
#400 value1=32'd71;value2=32'd78;
#400 value1=32'd81;value2=32'd84;
#400 value1=32'd91;value2=32'd94;
#400 value1=32'd96;value2=32'd102;
#400 value1=32'd103;value2=32'd183;
#400 value1=32'd261;value2=32'd382;
#400 value1=32'd427;value2=32'd512;
#400 value1=32'd25;value2=32'd44;
#400 value1=32'd63;value2=32'd82;
#400 value1=32'd90;value2=32'd91;
#400 value1=32'd94;value2=32'd97;
#400 value1=32'd104;value2=32'd184;
#400 value1=32'd262;value2=32'd383;
#400 value1=32'd428;value2=32'd513;
#400 value1=32'd26;value2=32'd54;
#400 value1=32'd71;value2=32'd83;
#400 value1=32'd90;value2=32'd92;
#400 value1=32'd93;value2=32'd98;
#400 value1=32'd104;value2=32'd185;
#400 value1=32'd263;value2=32'd384;
#400 value1=32'd429;value2=32'd514;
#400 value1=32'd10;value2=32'd35;
#400 value1=32'd45;value2=32'd64;
#400 value1=32'd79;value2=32'd85;
#400 value1=32'd86;value2=32'd91;
#400 value1=32'd96;value2=32'd97;
#400 value1=32'd100;value2=32'd101;
#400 value1=32'd186;value2=32'd264;
#400 value1=32'd385;value2=32'd430;
#400 value1=32'd515;value2=32'd540;
#400 value1=32'd11;value2=32'd36;
#400 value1=32'd55;value2=32'd72;
#400 value1=32'd79;value2=32'd85;
#400 value1=32'd87;value2=32'd92;
#400 value1=32'd95;value2=32'd98;
#400 value1=32'd102;value2=32'd103;
#400 value1=32'd187;value2=32'd265;
#400 value1=32'd386;value2=32'd431;
#400 value1=32'd516;value2=32'd541;
#400 value1=32'd12;value2=32'd37;
#400 value1=32'd45;value2=32'd64;
#400 value1=32'd88;value2=32'd90;
#400 value1=32'd93;value2=32'd95;
#400 value1=32'd98;value2=32'd104;
#400 value1=32'd188;value2=32'd266;
#400 value1=32'd387;value2=32'd432;
#400 value1=32'd517;value2=32'd542;
#400 value1=32'd13;value2=32'd38;
#400 value1=32'd55;value2=32'd72;
#400 value1=32'd89;value2=32'd90;
#400 value1=32'd94;value2=32'd96;
#400 value1=32'd97;value2=32'd104;
#400 value1=32'd189;value2=32'd267;
#400 value1=32'd388;value2=32'd433;
#400 value1=32'd518;value2=32'd543;
#400 value1=32'd47;value2=32'd56;
#400 value1=32'd66;value2=32'd73;
#400 value1=32'd80;value2=32'd81;
#400 value1=32'd86;value2=32'd87;
#400 value1=32'd101;value2=32'd102;
#400 value1=32'd190;value2=32'd268;
#400 value1=32'd389;value2=32'd434;
#400 value1=32'd519;value2=32'd544;
#400 value1=32'd46;value2=32'd48;
#400 value1=32'd65;value2=32'd67;
#400 value1=32'd82;value2=32'd88;
#400 value1=32'd91;value2=32'd95;
#400 value1=32'd101;value2=32'd102;
#400 value1=32'd191;value2=32'd269;
#400 value1=32'd390;value2=32'd435;
#400 value1=32'd520;value2=32'd545;
#400 value1=32'd49;value2=32'd56;
#400 value1=32'd68;value2=32'd73;
#400 value1=32'd83;value2=32'd89;
#400 value1=32'd91;value2=32'd95;
#400 value1=32'd99;value2=32'd100;
#400 value1=32'd103;value2=32'd104;
#400 value1=32'd192;value2=32'd270;
#400 value1=32'd391;value2=32'd436;
#400 value1=32'd521;value2=32'd546;
#400 value1=32'd47;value2=32'd58;
#400 value1=32'd66;value2=32'd75;
#400 value1=32'd82;value2=32'd88;
#400 value1=32'd92;value2=32'd96;
#400 value1=32'd99;value2=32'd100;
#400 value1=32'd103;value2=32'd104;
#400 value1=32'd193;value2=32'd271;
#400 value1=32'd392;value2=32'd437;
#400 value1=32'd522;value2=32'd547;
#400 value1=32'd57;value2=32'd59;
#400 value1=32'd74;value2=32'd76;
#400 value1=32'd83;value2=32'd89;
#400 value1=32'd92;value2=32'd96;
#400 value1=32'd101;value2=32'd102;
#400 value1=32'd194;value2=32'd272;
#400 value1=32'd393;value2=32'd438;
#400 value1=32'd523;value2=32'd548;
#400 value1=32'd49;value2=32'd58;
#400 value1=32'd68;value2=32'd75;
#400 value1=32'd93;value2=32'd94;
#400 value1=32'd97;value2=32'd98;
#400 value1=32'd101;value2=32'd102;
#400 value1=32'd195;value2=32'd273;
#400 value1=32'd394;value2=32'd439;
#400 value1=32'd524;value2=32'd549;
#400 value1=32'd1;value2=32'd14;
#400 value1=32'd108;value2=32'd109;
#400 value1=32'd111;value2=32'd113;
#400 value1=32'd120;value2=32'd121;
#400 value1=32'd122;value2=32'd124;
#400 value1=32'd196;value2=32'd197;
#400 value1=32'd201;value2=32'd203;
#400 value1=32'd0;value2=32'd2;
#400 value1=32'd15;value2=32'd107;
#400 value1=32'd108;value2=32'd114;
#400 value1=32'd116;value2=32'd118;
#400 value1=32'd131;value2=32'd132;
#400 value1=32'd133;value2=32'd135;
#400 value1=32'd196;value2=32'd208;
#400 value1=32'd212;value2=32'd214;
#400 value1=32'd0;value2=32'd3;
#400 value1=32'd16;value2=32'd106;
#400 value1=32'd109;value2=32'd115;
#400 value1=32'd117;value2=32'd119;
#400 value1=32'd141;value2=32'd142;
#400 value1=32'd143;value2=32'd145;
#400 value1=32'd197;value2=32'd208;
#400 value1=32'd222;value2=32'd224;
#400 value1=32'd4;value2=32'd17;
#400 value1=32'd105;value2=32'd106;
#400 value1=32'd109;value2=32'd114;
#400 value1=32'd116;value2=32'd120;
#400 value1=32'd151;value2=32'd152;
#400 value1=32'd154;value2=32'd198;
#400 value1=32'd209;value2=32'd219;
#400 value1=32'd231;value2=32'd233;
#400 value1=32'd5;value2=32'd18;
#400 value1=32'd105;value2=32'd107;
#400 value1=32'd108;value2=32'd115;
#400 value1=32'd117;value2=32'd121;
#400 value1=32'd151;value2=32'd160;
#400 value1=32'd162;value2=32'd199;
#400 value1=32'd210;value2=32'd220;
#400 value1=32'd239;value2=32'd241;
#400 value1=32'd0;value2=32'd6;
#400 value1=32'd19;value2=32'd111;
#400 value1=32'd112;value2=32'd114;
#400 value1=32'd115;value2=32'd122;
#400 value1=32'd152;value2=32'd160;
#400 value1=32'd169;value2=32'd200;
#400 value1=32'd211;value2=32'd221;
#400 value1=32'd246;value2=32'd248;
#400 value1=32'd7;value2=32'd20;
#400 value1=32'd105;value2=32'd110;
#400 value1=32'd113;value2=32'd114;
#400 value1=32'd115;value2=32'd123;
#400 value1=32'd153;value2=32'd161;
#400 value1=32'd168;value2=32'd175;
#400 value1=32'd201;value2=32'd212;
#400 value1=32'd222;value2=32'd254;
#400 value1=32'd0;value2=32'd8;
#400 value1=32'd21;value2=32'd110;
#400 value1=32'd113;value2=32'd116;
#400 value1=32'd117;value2=32'd124;
#400 value1=32'd154;value2=32'd162;
#400 value1=32'd169;value2=32'd202;
#400 value1=32'd213;value2=32'd223;
#400 value1=32'd253;value2=32'd259;
#400 value1=32'd9;value2=32'd22;
#400 value1=32'd105;value2=32'd111;
#400 value1=32'd112;value2=32'd116;
#400 value1=32'd117;value2=32'd125;
#400 value1=32'd155;value2=32'd163;
#400 value1=32'd170;value2=32'd181;
#400 value1=32'd203;value2=32'd214;
#400 value1=32'd224;value2=32'd254;
#400 value1=32'd10;value2=32'd23;
#400 value1=32'd106;value2=32'd108;
#400 value1=32'd110;value2=32'd111;
#400 value1=32'd115;value2=32'd116;
#400 value1=32'd126;value2=32'd156;
#400 value1=32'd164;value2=32'd171;
#400 value1=32'd182;value2=32'd204;
#400 value1=32'd215;value2=32'd225;
#400 value1=32'd255;value2=32'd264;
#400 value1=32'd11;value2=32'd24;
#400 value1=32'd107;value2=32'd109;
#400 value1=32'd110;value2=32'd111;
#400 value1=32'd114;value2=32'd117;
#400 value1=32'd127;value2=32'd157;
#400 value1=32'd165;value2=32'd172;
#400 value1=32'd183;value2=32'd205;
#400 value1=32'd216;value2=32'd226;
#400 value1=32'd256;value2=32'd265;
#400 value1=32'd12;value2=32'd25;
#400 value1=32'd106;value2=32'd108;
#400 value1=32'd112;value2=32'd113;
#400 value1=32'd114;value2=32'd117;
#400 value1=32'd128;value2=32'd158;
#400 value1=32'd166;value2=32'd173;
#400 value1=32'd184;value2=32'd206;
#400 value1=32'd217;value2=32'd227;
#400 value1=32'd257;value2=32'd266;
#400 value1=32'd13;value2=32'd26;
#400 value1=32'd107;value2=32'd109;
#400 value1=32'd112;value2=32'd113;
#400 value1=32'd115;value2=32'd116;
#400 value1=32'd129;value2=32'd159;
#400 value1=32'd167;value2=32'd174;
#400 value1=32'd185;value2=32'd207;
#400 value1=32'd218;value2=32'd228;
#400 value1=32'd258;value2=32'd267;
#400 value1=32'd1;value2=32'd27;
#400 value1=32'd106;value2=32'd119;
#400 value1=32'd120;value2=32'd126;
#400 value1=32'd128;value2=32'd131;
#400 value1=32'd132;value2=32'd134;
#400 value1=32'd136;value2=32'd274;
#400 value1=32'd278;value2=32'd280;
#400 value1=32'd1;value2=32'd28;
#400 value1=32'd107;value2=32'd118;
#400 value1=32'd121;value2=32'd127;
#400 value1=32'd129;value2=32'd141;
#400 value1=32'd142;value2=32'd144;
#400 value1=32'd146;value2=32'd274;
#400 value1=32'd288;value2=32'd290;
#400 value1=32'd29;value2=32'd105;
#400 value1=32'd108;value2=32'd118;
#400 value1=32'd121;value2=32'd126;
#400 value1=32'd128;value2=32'd151;
#400 value1=32'd153;value2=32'd155;
#400 value1=32'd275;value2=32'd285;
#400 value1=32'd297;value2=32'd299;
#400 value1=32'd30;value2=32'd105;
#400 value1=32'd109;value2=32'd119;
#400 value1=32'd120;value2=32'd127;
#400 value1=32'd129;value2=32'd151;
#400 value1=32'd161;value2=32'd163;
#400 value1=32'd276;value2=32'd286;
#400 value1=32'd305;value2=32'd307;
#400 value1=32'd1;value2=32'd31;
#400 value1=32'd105;value2=32'd110;
#400 value1=32'd123;value2=32'd124;
#400 value1=32'd126;value2=32'd127;
#400 value1=32'd152;value2=32'd160;
#400 value1=32'd168;value2=32'd170;
#400 value1=32'd277;value2=32'd287;
#400 value1=32'd312;value2=32'd314;
#400 value1=32'd32;value2=32'd111;
#400 value1=32'd122;value2=32'd125;
#400 value1=32'd126;value2=32'd127;
#400 value1=32'd153;value2=32'd161;
#400 value1=32'd176;value2=32'd278;
#400 value1=32'd288;value2=32'd320;
#400 value1=32'd1;value2=32'd33;
#400 value1=32'd105;value2=32'd112;
#400 value1=32'd122;value2=32'd125;
#400 value1=32'd128;value2=32'd129;
#400 value1=32'd154;value2=32'd162;
#400 value1=32'd175;value2=32'd181;
#400 value1=32'd279;value2=32'd289;
#400 value1=32'd319;value2=32'd325;
#400 value1=32'd34;value2=32'd113;
#400 value1=32'd123;value2=32'd124;
#400 value1=32'd128;value2=32'd129;
#400 value1=32'd155;value2=32'd163;
#400 value1=32'd176;value2=32'd280;
#400 value1=32'd290;value2=32'd320;
#400 value1=32'd35;value2=32'd114;
#400 value1=32'd118;value2=32'd120;
#400 value1=32'd122;value2=32'd123;
#400 value1=32'd127;value2=32'd128;
#400 value1=32'd156;value2=32'd164;
#400 value1=32'd177;value2=32'd186;
#400 value1=32'd281;value2=32'd291;
#400 value1=32'd321;value2=32'd330;
#400 value1=32'd36;value2=32'd115;
#400 value1=32'd119;value2=32'd121;
#400 value1=32'd122;value2=32'd123;
#400 value1=32'd126;value2=32'd129;
#400 value1=32'd157;value2=32'd165;
#400 value1=32'd178;value2=32'd187;
#400 value1=32'd282;value2=32'd292;
#400 value1=32'd322;value2=32'd331;
#400 value1=32'd37;value2=32'd116;
#400 value1=32'd118;value2=32'd120;
#400 value1=32'd124;value2=32'd125;
#400 value1=32'd126;value2=32'd129;
#400 value1=32'd158;value2=32'd166;
#400 value1=32'd179;value2=32'd188;
#400 value1=32'd283;value2=32'd293;
#400 value1=32'd323;value2=32'd332;
#400 value1=32'd38;value2=32'd117;
#400 value1=32'd119;value2=32'd121;
#400 value1=32'd124;value2=32'd125;
#400 value1=32'd127;value2=32'd128;
#400 value1=32'd159;value2=32'd167;
#400 value1=32'd180;value2=32'd189;
#400 value1=32'd284;value2=32'd294;
#400 value1=32'd324;value2=32'd333;
#400 value1=32'd2;value2=32'd3;
#400 value1=32'd39;value2=32'd132;
#400 value1=32'd138;value2=32'd140;
#400 value1=32'd141;value2=32'd147;
#400 value1=32'd149;value2=32'd274;
#400 value1=32'd343;value2=32'd345;
#400 value1=32'd4;value2=32'd40;
#400 value1=32'd106;value2=32'd118;
#400 value1=32'd132;value2=32'd137;
#400 value1=32'd139;value2=32'd141;
#400 value1=32'd156;value2=32'd158;
#400 value1=32'd275;value2=32'd340;
#400 value1=32'd352;value2=32'd354;
#400 value1=32'd5;value2=32'd41;
#400 value1=32'd106;value2=32'd118;
#400 value1=32'd130;value2=32'd131;
#400 value1=32'd138;value2=32'd140;
#400 value1=32'd142;value2=32'd151;
#400 value1=32'd164;value2=32'd166;
#400 value1=32'd276;value2=32'd341;
#400 value1=32'd360;value2=32'd362;
#400 value1=32'd2;value2=32'd6;
#400 value1=32'd42;value2=32'd106;
#400 value1=32'd134;value2=32'd135;
#400 value1=32'd137;value2=32'd138;
#400 value1=32'd143;value2=32'd152;
#400 value1=32'd171;value2=32'd173;
#400 value1=32'd277;value2=32'd342;
#400 value1=32'd367;value2=32'd369;
#400 value1=32'd7;value2=32'd43;
#400 value1=32'd118;value2=32'd133;
#400 value1=32'd136;value2=32'd137;
#400 value1=32'd138;value2=32'd144;
#400 value1=32'd153;value2=32'd177;
#400 value1=32'd179;value2=32'd278;
#400 value1=32'd343;value2=32'd375;
#400 value1=32'd2;value2=32'd8;
#400 value1=32'd44;value2=32'd106;
#400 value1=32'd133;value2=32'd136;
#400 value1=32'd139;value2=32'd140;
#400 value1=32'd145;value2=32'd154;
#400 value1=32'd182;value2=32'd184;
#400 value1=32'd279;value2=32'd344;
#400 value1=32'd374;value2=32'd380;
#400 value1=32'd9;value2=32'd45;
#400 value1=32'd118;value2=32'd134;
#400 value1=32'd135;value2=32'd139;
#400 value1=32'd140;value2=32'd146;
#400 value1=32'd155;value2=32'd186;
#400 value1=32'd188;value2=32'd280;
#400 value1=32'd345;value2=32'd375;
#400 value1=32'd10;value2=32'd46;
#400 value1=32'd131;value2=32'd133;
#400 value1=32'd134;value2=32'd138;
#400 value1=32'd139;value2=32'd147;
#400 value1=32'd156;value2=32'd191;
#400 value1=32'd281;value2=32'd346;
#400 value1=32'd376;value2=32'd385;
#400 value1=32'd11;value2=32'd47;
#400 value1=32'd130;value2=32'd132;
#400 value1=32'd133;value2=32'd134;
#400 value1=32'd137;value2=32'd140;
#400 value1=32'd148;value2=32'd157;
#400 value1=32'd190;value2=32'd193;
#400 value1=32'd282;value2=32'd347;
#400 value1=32'd377;value2=32'd386;
#400 value1=32'd12;value2=32'd48;
#400 value1=32'd131;value2=32'd135;
#400 value1=32'd136;value2=32'd137;
#400 value1=32'd140;value2=32'd149;
#400 value1=32'd158;value2=32'd191;
#400 value1=32'd283;value2=32'd348;
#400 value1=32'd378;value2=32'd387;
#400 value1=32'd13;value2=32'd49;
#400 value1=32'd130;value2=32'd132;
#400 value1=32'd135;value2=32'd136;
#400 value1=32'd138;value2=32'd139;
#400 value1=32'd150;value2=32'd159;
#400 value1=32'd192;value2=32'd195;
#400 value1=32'd284;value2=32'd349;
#400 value1=32'd379;value2=32'd388;
#400 value1=32'd4;value2=32'd50;
#400 value1=32'd107;value2=32'd119;
#400 value1=32'd130;value2=32'd131;
#400 value1=32'd142;value2=32'd147;
#400 value1=32'd149;value2=32'd151;
#400 value1=32'd157;value2=32'd159;
#400 value1=32'd285;value2=32'd340;
#400 value1=32'd397;value2=32'd399;
#400 value1=32'd5;value2=32'd51;
#400 value1=32'd107;value2=32'd119;
#400 value1=32'd132;value2=32'd141;
#400 value1=32'd148;value2=32'd150;
#400 value1=32'd165;value2=32'd167;
#400 value1=32'd286;value2=32'd341;
#400 value1=32'd405;value2=32'd407;
#400 value1=32'd3;value2=32'd6;
#400 value1=32'd52;value2=32'd107;
#400 value1=32'd133;value2=32'd144;
#400 value1=32'd145;value2=32'd147;
#400 value1=32'd148;value2=32'd160;
#400 value1=32'd172;value2=32'd174;
#400 value1=32'd287;value2=32'd342;
#400 value1=32'd412;value2=32'd414;
#400 value1=32'd7;value2=32'd53;
#400 value1=32'd119;value2=32'd134;
#400 value1=32'd143;value2=32'd146;
#400 value1=32'd147;value2=32'd148;
#400 value1=32'd161;value2=32'd178;
#400 value1=32'd180;value2=32'd288;
#400 value1=32'd343;value2=32'd420;
#400 value1=32'd3;value2=32'd8;
#400 value1=32'd54;value2=32'd107;
#400 value1=32'd135;value2=32'd143;
#400 value1=32'd146;value2=32'd149;
#400 value1=32'd150;value2=32'd162;
#400 value1=32'd183;value2=32'd185;
#400 value1=32'd289;value2=32'd344;
#400 value1=32'd419;value2=32'd425;
#400 value1=32'd9;value2=32'd55;
#400 value1=32'd119;value2=32'd136;
#400 value1=32'd144;value2=32'd145;
#400 value1=32'd149;value2=32'd150;
#400 value1=32'd163;value2=32'd187;
#400 value1=32'd189;value2=32'd290;
#400 value1=32'd345;value2=32'd420;
#400 value1=32'd10;value2=32'd56;
#400 value1=32'd130;value2=32'd137;
#400 value1=32'd141;value2=32'd143;
#400 value1=32'd144;value2=32'd148;
#400 value1=32'd149;value2=32'd164;
#400 value1=32'd190;value2=32'd192;
#400 value1=32'd291;value2=32'd346;
#400 value1=32'd421;value2=32'd430;
#400 value1=32'd11;value2=32'd57;
#400 value1=32'd138;value2=32'd142;
#400 value1=32'd143;value2=32'd144;
#400 value1=32'd147;value2=32'd150;
#400 value1=32'd165;value2=32'd194;
#400 value1=32'd292;value2=32'd347;
#400 value1=32'd422;value2=32'd431;
#400 value1=32'd12;value2=32'd58;
#400 value1=32'd130;value2=32'd139;
#400 value1=32'd141;value2=32'd145;
#400 value1=32'd146;value2=32'd147;
#400 value1=32'd150;value2=32'd166;
#400 value1=32'd193;value2=32'd195;
#400 value1=32'd293;value2=32'd348;
#400 value1=32'd423;value2=32'd432;
#400 value1=32'd13;value2=32'd59;
#400 value1=32'd140;value2=32'd142;
#400 value1=32'd145;value2=32'd146;
#400 value1=32'd148;value2=32'd149;
#400 value1=32'd167;value2=32'd194;
#400 value1=32'd294;value2=32'd349;
#400 value1=32'd424;value2=32'd433;
#400 value1=32'd60;value2=32'd108;
#400 value1=32'd109;value2=32'd120;
#400 value1=32'd121;value2=32'd132;
#400 value1=32'd141;value2=32'd157;
#400 value1=32'd159;value2=32'd164;
#400 value1=32'd166;value2=32'd295;
#400 value1=32'd350;value2=32'd395;
#400 value1=32'd441;value2=32'd443;
#400 value1=32'd4;value2=32'd61;
#400 value1=32'd108;value2=32'd110;
#400 value1=32'd122;value2=32'd133;
#400 value1=32'd153;value2=32'd154;
#400 value1=32'd156;value2=32'd157;
#400 value1=32'd160;value2=32'd171;
#400 value1=32'd173;value2=32'd296;
#400 value1=32'd351;value2=32'd396;
#400 value1=32'd448;value2=32'd450;
#400 value1=32'd62;value2=32'd111;
#400 value1=32'd120;value2=32'd123;
#400 value1=32'd134;value2=32'd152;
#400 value1=32'd155;value2=32'd156;
#400 value1=32'd157;value2=32'd161;
#400 value1=32'd177;value2=32'd179;
#400 value1=32'd297;value2=32'd352;
#400 value1=32'd397;value2=32'd456;
#400 value1=32'd4;value2=32'd63;
#400 value1=32'd108;value2=32'd112;
#400 value1=32'd124;value2=32'd135;
#400 value1=32'd152;value2=32'd155;
#400 value1=32'd158;value2=32'd159;
#400 value1=32'd162;value2=32'd182;
#400 value1=32'd184;value2=32'd298;
#400 value1=32'd353;value2=32'd398;
#400 value1=32'd455;value2=32'd461;
#400 value1=32'd64;value2=32'd113;
#400 value1=32'd120;value2=32'd125;
#400 value1=32'd136;value2=32'd153;
#400 value1=32'd154;value2=32'd158;
#400 value1=32'd159;value2=32'd163;
#400 value1=32'd186;value2=32'd188;
#400 value1=32'd299;value2=32'd354;
#400 value1=32'd399;value2=32'd456;
#400 value1=32'd65;value2=32'd114;
#400 value1=32'd126;value2=32'd131;
#400 value1=32'd137;value2=32'd152;
#400 value1=32'd153;value2=32'd157;
#400 value1=32'd158;value2=32'd164;
#400 value1=32'd191;value2=32'd300;
#400 value1=32'd355;value2=32'd400;
#400 value1=32'd457;value2=32'd466;
#400 value1=32'd66;value2=32'd115;
#400 value1=32'd127;value2=32'd138;
#400 value1=32'd141;value2=32'd151;
#400 value1=32'd152;value2=32'd153;
#400 value1=32'd156;value2=32'd159;
#400 value1=32'd165;value2=32'd190;
#400 value1=32'd193;value2=32'd301;
#400 value1=32'd356;value2=32'd401;
#400 value1=32'd458;value2=32'd467;
#400 value1=32'd67;value2=32'd116;
#400 value1=32'd128;value2=32'd131;
#400 value1=32'd139;value2=32'd154;
#400 value1=32'd155;value2=32'd156;
#400 value1=32'd159;value2=32'd166;
#400 value1=32'd191;value2=32'd302;
#400 value1=32'd357;value2=32'd402;
#400 value1=32'd459;value2=32'd468;
#400 value1=32'd68;value2=32'd117;
#400 value1=32'd129;value2=32'd140;
#400 value1=32'd141;value2=32'd151;
#400 value1=32'd154;value2=32'd155;
#400 value1=32'd157;value2=32'd158;
#400 value1=32'd167;value2=32'd192;
#400 value1=32'd195;value2=32'd303;
#400 value1=32'd358;value2=32'd403;
#400 value1=32'd460;value2=32'd469;
#400 value1=32'd5;value2=32'd69;
#400 value1=32'd109;value2=32'd110;
#400 value1=32'd122;value2=32'd143;
#400 value1=32'd152;value2=32'd161;
#400 value1=32'd162;value2=32'd164;
#400 value1=32'd165;value2=32'd172;
#400 value1=32'd174;value2=32'd304;
#400 value1=32'd359;value2=32'd404;
#400 value1=32'd476;value2=32'd478;
#400 value1=32'd70;value2=32'd111;
#400 value1=32'd121;value2=32'd123;
#400 value1=32'd144;value2=32'd153;
#400 value1=32'd160;value2=32'd163;
#400 value1=32'd164;value2=32'd165;
#400 value1=32'd178;value2=32'd180;
#400 value1=32'd305;value2=32'd360;
#400 value1=32'd405;value2=32'd484;
#400 value1=32'd5;value2=32'd71;
#400 value1=32'd109;value2=32'd112;
#400 value1=32'd124;value2=32'd145;
#400 value1=32'd154;value2=32'd160;
#400 value1=32'd163;value2=32'd166;
#400 value1=32'd167;value2=32'd183;
#400 value1=32'd185;value2=32'd306;
#400 value1=32'd361;value2=32'd406;
#400 value1=32'd483;value2=32'd489;
#400 value1=32'd72;value2=32'd113;
#400 value1=32'd121;value2=32'd125;
#400 value1=32'd146;value2=32'd155;
#400 value1=32'd161;value2=32'd162;
#400 value1=32'd166;value2=32'd167;
#400 value1=32'd187;value2=32'd189;
#400 value1=32'd307;value2=32'd362;
#400 value1=32'd407;value2=32'd484;
#400 value1=32'd73;value2=32'd114;
#400 value1=32'd126;value2=32'd132;
#400 value1=32'd147;value2=32'd151;
#400 value1=32'd156;value2=32'd160;
#400 value1=32'd161;value2=32'd165;
#400 value1=32'd166;value2=32'd190;
#400 value1=32'd192;value2=32'd308;
#400 value1=32'd363;value2=32'd408;
#400 value1=32'd485;value2=32'd494;
#400 value1=32'd74;value2=32'd115;
#400 value1=32'd127;value2=32'd142;
#400 value1=32'd148;value2=32'd157;
#400 value1=32'd160;value2=32'd161;
#400 value1=32'd164;value2=32'd167;
#400 value1=32'd194;value2=32'd309;
#400 value1=32'd364;value2=32'd409;
#400 value1=32'd486;value2=32'd495;
#400 value1=32'd75;value2=32'd116;
#400 value1=32'd128;value2=32'd132;
#400 value1=32'd149;value2=32'd151;
#400 value1=32'd158;value2=32'd162;
#400 value1=32'd163;value2=32'd164;
#400 value1=32'd167;value2=32'd193;
#400 value1=32'd195;value2=32'd310;
#400 value1=32'd365;value2=32'd410;
#400 value1=32'd487;value2=32'd496;
#400 value1=32'd76;value2=32'd117;
#400 value1=32'd129;value2=32'd142;
#400 value1=32'd150;value2=32'd159;
#400 value1=32'd162;value2=32'd163;
#400 value1=32'd165;value2=32'd166;
#400 value1=32'd194;value2=32'd311;
#400 value1=32'd366;value2=32'd411;
#400 value1=32'd488;value2=32'd497;
#400 value1=32'd7;value2=32'd77;
#400 value1=32'd111;value2=32'd122;
#400 value1=32'd170;value2=32'd171;
#400 value1=32'd172;value2=32'd175;
#400 value1=32'd177;value2=32'd178;
#400 value1=32'd312;value2=32'd367;
#400 value1=32'd412;value2=32'd505;
#400 value1=32'd6;value2=32'd8;
#400 value1=32'd78;value2=32'd110;
#400 value1=32'd112;value2=32'd170;
#400 value1=32'd173;value2=32'd174;
#400 value1=32'd175;value2=32'd182;
#400 value1=32'd183;value2=32'd313;
#400 value1=32'd368;value2=32'd413;
#400 value1=32'd504;value2=32'd510;
#400 value1=32'd9;value2=32'd79;
#400 value1=32'd113;value2=32'd122;
#400 value1=32'd168;value2=32'd169;
#400 value1=32'd173;value2=32'd174;
#400 value1=32'd176;value2=32'd181;
#400 value1=32'd186;value2=32'd187;
#400 value1=32'd314;value2=32'd369;
#400 value1=32'd414;value2=32'd505;
#400 value1=32'd10;value2=32'd80;
#400 value1=32'd114;value2=32'd133;
#400 value1=32'd152;value2=32'd168;
#400 value1=32'd172;value2=32'd173;
#400 value1=32'd177;value2=32'd182;
#400 value1=32'd190;value2=32'd315;
#400 value1=32'd370;value2=32'd415;
#400 value1=32'd506;value2=32'd515;
#400 value1=32'd11;value2=32'd81;
#400 value1=32'd115;value2=32'd143;
#400 value1=32'd160;value2=32'd168;
#400 value1=32'd171;value2=32'd174;
#400 value1=32'd178;value2=32'd183;
#400 value1=32'd190;value2=32'd316;
#400 value1=32'd371;value2=32'd416;
#400 value1=32'd507;value2=32'd516;
#400 value1=32'd12;value2=32'd82;
#400 value1=32'd116;value2=32'd133;
#400 value1=32'd152;value2=32'd169;
#400 value1=32'd170;value2=32'd171;
#400 value1=32'd174;value2=32'd179;
#400 value1=32'd184;value2=32'd191;
#400 value1=32'd193;value2=32'd317;
#400 value1=32'd372;value2=32'd417;
#400 value1=32'd508;value2=32'd517;
#400 value1=32'd13;value2=32'd83;
#400 value1=32'd117;value2=32'd143;
#400 value1=32'd160;value2=32'd169;
#400 value1=32'd170;value2=32'd172;
#400 value1=32'd173;value2=32'd180;
#400 value1=32'd185;value2=32'd192;
#400 value1=32'd194;value2=32'd318;
#400 value1=32'd373;value2=32'd418;
#400 value1=32'd509;value2=32'd518;
#400 value1=32'd7;value2=32'd84;
#400 value1=32'd111;value2=32'd124;
#400 value1=32'd168;value2=32'd169;
#400 value1=32'd176;value2=32'd179;
#400 value1=32'd180;value2=32'd181;
#400 value1=32'd182;value2=32'd183;
#400 value1=32'd319;value2=32'd374;
#400 value1=32'd419;value2=32'd525;
#400 value1=32'd85;value2=32'd123;
#400 value1=32'd125;value2=32'd170;
#400 value1=32'd175;value2=32'd179;
#400 value1=32'd180;value2=32'd186;
#400 value1=32'd187;value2=32'd320;
#400 value1=32'd375;value2=32'd420;
#400 value1=32'd86;value2=32'd126;
#400 value1=32'd134;value2=32'd153;
#400 value1=32'd168;value2=32'd171;
#400 value1=32'd178;value2=32'd179;
#400 value1=32'd186;value2=32'd190;
#400 value1=32'd321;value2=32'd376;
#400 value1=32'd421;value2=32'd530;
#400 value1=32'd87;value2=32'd127;
#400 value1=32'd144;value2=32'd161;
#400 value1=32'd168;value2=32'd172;
#400 value1=32'd177;value2=32'd180;
#400 value1=32'd187;value2=32'd190;
#400 value1=32'd322;value2=32'd377;
#400 value1=32'd422;value2=32'd531;
#400 value1=32'd88;value2=32'd128;
#400 value1=32'd134;value2=32'd153;
#400 value1=32'd173;value2=32'd175;
#400 value1=32'd176;value2=32'd177;
#400 value1=32'd180;value2=32'd188;
#400 value1=32'd191;value2=32'd193;
#400 value1=32'd323;value2=32'd378;
#400 value1=32'd423;value2=32'd532;
#400 value1=32'd89;value2=32'd129;
#400 value1=32'd144;value2=32'd161;
#400 value1=32'd174;value2=32'd175;
#400 value1=32'd176;value2=32'd178;
#400 value1=32'd179;value2=32'd189;
#400 value1=32'd192;value2=32'd194;
#400 value1=32'd324;value2=32'd379;
#400 value1=32'd424;value2=32'd533;
#400 value1=32'd9;value2=32'd90;
#400 value1=32'd113;value2=32'd124;
#400 value1=32'd170;value2=32'd175;
#400 value1=32'd184;value2=32'd185;
#400 value1=32'd188;value2=32'd189;
#400 value1=32'd325;value2=32'd380;
#400 value1=32'd425;value2=32'd525;
#400 value1=32'd10;value2=32'd91;
#400 value1=32'd114;value2=32'd135;
#400 value1=32'd154;value2=32'd169;
#400 value1=32'd171;value2=32'd175;
#400 value1=32'd183;value2=32'd184;
#400 value1=32'd186;value2=32'd191;
#400 value1=32'd192;value2=32'd326;
#400 value1=32'd381;value2=32'd426;
#400 value1=32'd526;value2=32'd540;
#400 value1=32'd11;value2=32'd92;
#400 value1=32'd115;value2=32'd145;
#400 value1=32'd162;value2=32'd169;
#400 value1=32'd172;value2=32'd175;
#400 value1=32'd182;value2=32'd185;
#400 value1=32'd187;value2=32'd193;
#400 value1=32'd194;value2=32'd327;
#400 value1=32'd382;value2=32'd427;
#400 value1=32'd527;value2=32'd541;
#400 value1=32'd12;value2=32'd93;
#400 value1=32'd116;value2=32'd135;
#400 value1=32'd154;value2=32'd173;
#400 value1=32'd181;value2=32'd182;
#400 value1=32'd185;value2=32'd188;
#400 value1=32'd195;value2=32'd328;
#400 value1=32'd383;value2=32'd428;
#400 value1=32'd528;value2=32'd542;
#400 value1=32'd13;value2=32'd94;
#400 value1=32'd117;value2=32'd145;
#400 value1=32'd162;value2=32'd174;
#400 value1=32'd181;value2=32'd183;
#400 value1=32'd184;value2=32'd189;
#400 value1=32'd195;value2=32'd329;
#400 value1=32'd384;value2=32'd429;
#400 value1=32'd529;value2=32'd543;
#400 value1=32'd95;value2=32'd126;
#400 value1=32'd136;value2=32'd155;
#400 value1=32'd170;value2=32'd176;
#400 value1=32'd177;value2=32'd182;
#400 value1=32'd187;value2=32'd188;
#400 value1=32'd191;value2=32'd192;
#400 value1=32'd330;value2=32'd385;
#400 value1=32'd430;value2=32'd530;
#400 value1=32'd96;value2=32'd127;
#400 value1=32'd146;value2=32'd163;
#400 value1=32'd170;value2=32'd176;
#400 value1=32'd178;value2=32'd183;
#400 value1=32'd186;value2=32'd189;
#400 value1=32'd193;value2=32'd194;
#400 value1=32'd331;value2=32'd386;
#400 value1=32'd431;value2=32'd531;
#400 value1=32'd97;value2=32'd128;
#400 value1=32'd136;value2=32'd155;
#400 value1=32'd179;value2=32'd181;
#400 value1=32'd184;value2=32'd186;
#400 value1=32'd189;value2=32'd195;
#400 value1=32'd332;value2=32'd387;
#400 value1=32'd432;value2=32'd532;
#400 value1=32'd98;value2=32'd129;
#400 value1=32'd146;value2=32'd163;
#400 value1=32'd180;value2=32'd181;
#400 value1=32'd185;value2=32'd187;
#400 value1=32'd188;value2=32'd195;
#400 value1=32'd333;value2=32'd388;
#400 value1=32'd433;value2=32'd533;
#400 value1=32'd99;value2=32'd138;
#400 value1=32'd147;value2=32'd157;
#400 value1=32'd164;value2=32'd171;
#400 value1=32'd172;value2=32'd177;
#400 value1=32'd178;value2=32'd192;
#400 value1=32'd193;value2=32'd334;
#400 value1=32'd389;value2=32'd434;
#400 value1=32'd534;value2=32'd550;
#400 value1=32'd100;value2=32'd137;
#400 value1=32'd139;value2=32'd156;
#400 value1=32'd158;value2=32'd173;
#400 value1=32'd179;value2=32'd182;
#400 value1=32'd186;value2=32'd192;
#400 value1=32'd193;value2=32'd335;
#400 value1=32'd390;value2=32'd435;
#400 value1=32'd535;value2=32'd551;
#400 value1=32'd101;value2=32'd140;
#400 value1=32'd147;value2=32'd159;
#400 value1=32'd164;value2=32'd174;
#400 value1=32'd180;value2=32'd182;
#400 value1=32'd186;value2=32'd190;
#400 value1=32'd191;value2=32'd194;
#400 value1=32'd195;value2=32'd336;
#400 value1=32'd391;value2=32'd436;
#400 value1=32'd536;value2=32'd552;
#400 value1=32'd102;value2=32'd138;
#400 value1=32'd149;value2=32'd157;
#400 value1=32'd166;value2=32'd173;
#400 value1=32'd179;value2=32'd183;
#400 value1=32'd187;value2=32'd190;
#400 value1=32'd191;value2=32'd194;
#400 value1=32'd195;value2=32'd337;
#400 value1=32'd392;value2=32'd437;
#400 value1=32'd537;value2=32'd553;
#400 value1=32'd103;value2=32'd148;
#400 value1=32'd150;value2=32'd165;
#400 value1=32'd167;value2=32'd174;
#400 value1=32'd180;value2=32'd183;
#400 value1=32'd187;value2=32'd192;
#400 value1=32'd193;value2=32'd338;
#400 value1=32'd393;value2=32'd438;
#400 value1=32'd538;value2=32'd554;
#400 value1=32'd104;value2=32'd140;
#400 value1=32'd149;value2=32'd159;
#400 value1=32'd166;value2=32'd184;
#400 value1=32'd185;value2=32'd188;
#400 value1=32'd189;value2=32'd192;
#400 value1=32'd193;value2=32'd339;
#400 value1=32'd394;value2=32'd439;
#400 value1=32'd539;value2=32'd555;
#400 value1=32'd14;value2=32'd27;
#400 value1=32'd105;value2=32'd106;
#400 value1=32'd197;value2=32'd198;
#400 value1=32'd204;value2=32'd206;
#400 value1=32'd209;value2=32'd210;
#400 value1=32'd212;value2=32'd214;
#400 value1=32'd275;value2=32'd276;
#400 value1=32'd277;value2=32'd279;
#400 value1=32'd14;value2=32'd28;
#400 value1=32'd105;value2=32'd107;
#400 value1=32'd196;value2=32'd199;
#400 value1=32'd205;value2=32'd207;
#400 value1=32'd219;value2=32'd220;
#400 value1=32'd222;value2=32'd224;
#400 value1=32'd285;value2=32'd286;
#400 value1=32'd287;value2=32'd289;
#400 value1=32'd29;value2=32'd108;
#400 value1=32'd196;value2=32'd199;
#400 value1=32'd204;value2=32'd206;
#400 value1=32'd229;value2=32'd231;
#400 value1=32'd233;value2=32'd295;
#400 value1=32'd296;value2=32'd298;
#400 value1=32'd30;value2=32'd109;
#400 value1=32'd197;value2=32'd198;
#400 value1=32'd205;value2=32'd207;
#400 value1=32'd229;value2=32'd239;
#400 value1=32'd241;value2=32'd295;
#400 value1=32'd304;value2=32'd306;
#400 value1=32'd14;value2=32'd31;
#400 value1=32'd110;value2=32'd201;
#400 value1=32'd202;value2=32'd204;
#400 value1=32'd205;value2=32'd230;
#400 value1=32'd238;value2=32'd246;
#400 value1=32'd248;value2=32'd296;
#400 value1=32'd304;value2=32'd313;
#400 value1=32'd32;value2=32'd105;
#400 value1=32'd111;value2=32'd200;
#400 value1=32'd203;value2=32'd204;
#400 value1=32'd205;value2=32'd231;
#400 value1=32'd239;value2=32'd254;
#400 value1=32'd297;value2=32'd305;
#400 value1=32'd312;value2=32'd319;
#400 value1=32'd14;value2=32'd33;
#400 value1=32'd112;value2=32'd200;
#400 value1=32'd203;value2=32'd206;
#400 value1=32'd207;value2=32'd232;
#400 value1=32'd240;value2=32'd253;
#400 value1=32'd259;value2=32'd298;
#400 value1=32'd306;value2=32'd313;
#400 value1=32'd34;value2=32'd105;
#400 value1=32'd113;value2=32'd201;
#400 value1=32'd202;value2=32'd206;
#400 value1=32'd207;value2=32'd233;
#400 value1=32'd241;value2=32'd254;
#400 value1=32'd299;value2=32'd307;
#400 value1=32'd314;value2=32'd325;
#400 value1=32'd35;value2=32'd114;
#400 value1=32'd196;value2=32'd198;
#400 value1=32'd200;value2=32'd201;
#400 value1=32'd205;value2=32'd206;
#400 value1=32'd234;value2=32'd242;
#400 value1=32'd255;value2=32'd264;
#400 value1=32'd300;value2=32'd308;
#400 value1=32'd315;value2=32'd326;
#400 value1=32'd36;value2=32'd115;
#400 value1=32'd197;value2=32'd199;
#400 value1=32'd200;value2=32'd201;
#400 value1=32'd204;value2=32'd207;
#400 value1=32'd235;value2=32'd243;
#400 value1=32'd256;value2=32'd265;
#400 value1=32'd301;value2=32'd309;
#400 value1=32'd316;value2=32'd327;
#400 value1=32'd37;value2=32'd116;
#400 value1=32'd196;value2=32'd198;
#400 value1=32'd202;value2=32'd203;
#400 value1=32'd204;value2=32'd207;
#400 value1=32'd236;value2=32'd244;
#400 value1=32'd257;value2=32'd266;
#400 value1=32'd302;value2=32'd310;
#400 value1=32'd317;value2=32'd328;
#400 value1=32'd38;value2=32'd117;
#400 value1=32'd197;value2=32'd199;
#400 value1=32'd202;value2=32'd203;
#400 value1=32'd205;value2=32'd206;
#400 value1=32'd237;value2=32'd245;
#400 value1=32'd258;value2=32'd267;
#400 value1=32'd303;value2=32'd311;
#400 value1=32'd318;value2=32'd329;
#400 value1=32'd15;value2=32'd16;
#400 value1=32'd39;value2=32'd106;
#400 value1=32'd107;value2=32'd210;
#400 value1=32'd216;value2=32'd218;
#400 value1=32'd219;value2=32'd225;
#400 value1=32'd227;value2=32'd274;
#400 value1=32'd340;value2=32'd341;
#400 value1=32'd342;value2=32'd344;
#400 value1=32'd17;value2=32'd40;
#400 value1=32'd108;value2=32'd196;
#400 value1=32'd210;value2=32'd215;
#400 value1=32'd217;value2=32'd219;
#400 value1=32'd234;value2=32'd236;
#400 value1=32'd275;value2=32'd350;
#400 value1=32'd351;value2=32'd353;
#400 value1=32'd18;value2=32'd41;
#400 value1=32'd109;value2=32'd196;
#400 value1=32'd208;value2=32'd209;
#400 value1=32'd216;value2=32'd218;
#400 value1=32'd220;value2=32'd229;
#400 value1=32'd242;value2=32'd244;
#400 value1=32'd276;value2=32'd350;
#400 value1=32'd359;value2=32'd361;
#400 value1=32'd15;value2=32'd19;
#400 value1=32'd42;value2=32'd110;
#400 value1=32'd212;value2=32'd213;
#400 value1=32'd215;value2=32'd216;
#400 value1=32'd221;value2=32'd230;
#400 value1=32'd249;value2=32'd251;
#400 value1=32'd277;value2=32'd351;
#400 value1=32'd359;value2=32'd368;
#400 value1=32'd20;value2=32'd43;
#400 value1=32'd106;value2=32'd111;
#400 value1=32'd196;value2=32'd211;
#400 value1=32'd214;value2=32'd215;
#400 value1=32'd216;value2=32'd222;
#400 value1=32'd231;value2=32'd255;
#400 value1=32'd257;value2=32'd278;
#400 value1=32'd352;value2=32'd360;
#400 value1=32'd367;value2=32'd374;
#400 value1=32'd15;value2=32'd21;
#400 value1=32'd44;value2=32'd112;
#400 value1=32'd211;value2=32'd214;
#400 value1=32'd217;value2=32'd218;
#400 value1=32'd223;value2=32'd232;
#400 value1=32'd260;value2=32'd262;
#400 value1=32'd279;value2=32'd353;
#400 value1=32'd361;value2=32'd368;
#400 value1=32'd22;value2=32'd45;
#400 value1=32'd106;value2=32'd113;
#400 value1=32'd196;value2=32'd212;
#400 value1=32'd213;value2=32'd217;
#400 value1=32'd218;value2=32'd224;
#400 value1=32'd233;value2=32'd264;
#400 value1=32'd266;value2=32'd280;
#400 value1=32'd354;value2=32'd362;
#400 value1=32'd369;value2=32'd380;
#400 value1=32'd23;value2=32'd46;
#400 value1=32'd114;value2=32'd209;
#400 value1=32'd211;value2=32'd212;
#400 value1=32'd216;value2=32'd217;
#400 value1=32'd225;value2=32'd234;
#400 value1=32'd269;value2=32'd281;
#400 value1=32'd355;value2=32'd363;
#400 value1=32'd370;value2=32'd381;
#400 value1=32'd24;value2=32'd47;
#400 value1=32'd115;value2=32'd208;
#400 value1=32'd210;value2=32'd211;
#400 value1=32'd212;value2=32'd215;
#400 value1=32'd218;value2=32'd226;
#400 value1=32'd235;value2=32'd268;
#400 value1=32'd271;value2=32'd282;
#400 value1=32'd356;value2=32'd364;
#400 value1=32'd371;value2=32'd382;
#400 value1=32'd25;value2=32'd48;
#400 value1=32'd116;value2=32'd209;
#400 value1=32'd213;value2=32'd214;
#400 value1=32'd215;value2=32'd218;
#400 value1=32'd227;value2=32'd236;
#400 value1=32'd269;value2=32'd283;
#400 value1=32'd357;value2=32'd365;
#400 value1=32'd372;value2=32'd383;
#400 value1=32'd26;value2=32'd49;
#400 value1=32'd117;value2=32'd208;
#400 value1=32'd210;value2=32'd213;
#400 value1=32'd214;value2=32'd216;
#400 value1=32'd217;value2=32'd228;
#400 value1=32'd237;value2=32'd270;
#400 value1=32'd273;value2=32'd284;
#400 value1=32'd358;value2=32'd366;
#400 value1=32'd373;value2=32'd384;
#400 value1=32'd17;value2=32'd50;
#400 value1=32'd108;value2=32'd197;
#400 value1=32'd208;value2=32'd209;
#400 value1=32'd220;value2=32'd225;
#400 value1=32'd227;value2=32'd229;
#400 value1=32'd235;value2=32'd237;
#400 value1=32'd285;value2=32'd395;
#400 value1=32'd396;value2=32'd398;
#400 value1=32'd18;value2=32'd51;
#400 value1=32'd109;value2=32'd197;
#400 value1=32'd210;value2=32'd219;
#400 value1=32'd226;value2=32'd228;
#400 value1=32'd243;value2=32'd245;
#400 value1=32'd286;value2=32'd395;
#400 value1=32'd404;value2=32'd406;
#400 value1=32'd16;value2=32'd19;
#400 value1=32'd52;value2=32'd110;
#400 value1=32'd211;value2=32'd222;
#400 value1=32'd223;value2=32'd225;
#400 value1=32'd226;value2=32'd238;
#400 value1=32'd250;value2=32'd252;
#400 value1=32'd287;value2=32'd396;
#400 value1=32'd404;value2=32'd413;
#400 value1=32'd20;value2=32'd53;
#400 value1=32'd107;value2=32'd111;
#400 value1=32'd197;value2=32'd212;
#400 value1=32'd221;value2=32'd224;
#400 value1=32'd225;value2=32'd226;
#400 value1=32'd239;value2=32'd256;
#400 value1=32'd258;value2=32'd288;
#400 value1=32'd397;value2=32'd405;
#400 value1=32'd412;value2=32'd419;
#400 value1=32'd16;value2=32'd21;
#400 value1=32'd54;value2=32'd112;
#400 value1=32'd213;value2=32'd221;
#400 value1=32'd224;value2=32'd227;
#400 value1=32'd228;value2=32'd240;
#400 value1=32'd261;value2=32'd263;
#400 value1=32'd289;value2=32'd398;
#400 value1=32'd406;value2=32'd413;
#400 value1=32'd22;value2=32'd55;
#400 value1=32'd107;value2=32'd113;
#400 value1=32'd197;value2=32'd214;
#400 value1=32'd222;value2=32'd223;
#400 value1=32'd227;value2=32'd228;
#400 value1=32'd241;value2=32'd265;
#400 value1=32'd267;value2=32'd290;
#400 value1=32'd399;value2=32'd407;
#400 value1=32'd414;value2=32'd425;
#400 value1=32'd23;value2=32'd56;
#400 value1=32'd114;value2=32'd208;
#400 value1=32'd215;value2=32'd219;
#400 value1=32'd221;value2=32'd222;
#400 value1=32'd226;value2=32'd227;
#400 value1=32'd242;value2=32'd268;
#400 value1=32'd270;value2=32'd291;
#400 value1=32'd400;value2=32'd408;
#400 value1=32'd415;value2=32'd426;
#400 value1=32'd24;value2=32'd57;
#400 value1=32'd115;value2=32'd216;
#400 value1=32'd220;value2=32'd221;
#400 value1=32'd222;value2=32'd225;
#400 value1=32'd228;value2=32'd243;
#400 value1=32'd272;value2=32'd292;
#400 value1=32'd401;value2=32'd409;
#400 value1=32'd416;value2=32'd427;
#400 value1=32'd25;value2=32'd58;
#400 value1=32'd116;value2=32'd208;
#400 value1=32'd217;value2=32'd219;
#400 value1=32'd223;value2=32'd224;
#400 value1=32'd225;value2=32'd228;
#400 value1=32'd244;value2=32'd271;
#400 value1=32'd273;value2=32'd293;
#400 value1=32'd402;value2=32'd410;
#400 value1=32'd417;value2=32'd428;
#400 value1=32'd26;value2=32'd59;
#400 value1=32'd117;value2=32'd218;
#400 value1=32'd220;value2=32'd223;
#400 value1=32'd224;value2=32'd226;
#400 value1=32'd227;value2=32'd245;
#400 value1=32'd272;value2=32'd294;
#400 value1=32'd403;value2=32'd411;
#400 value1=32'd418;value2=32'd429;
#400 value1=32'd60;value2=32'd198;
#400 value1=32'd199;value2=32'd210;
#400 value1=32'd219;value2=32'd235;
#400 value1=32'd237;value2=32'd242;
#400 value1=32'd244;value2=32'd295;
#400 value1=32'd440;value2=32'd442;
#400 value1=32'd17;value2=32'd61;
#400 value1=32'd200;value2=32'd211;
#400 value1=32'd231;value2=32'd232;
#400 value1=32'd234;value2=32'd235;
#400 value1=32'd238;value2=32'd249;
#400 value1=32'd251;value2=32'd296;
#400 value1=32'd440;value2=32'd449;
#400 value1=32'd62;value2=32'd108;
#400 value1=32'd198;value2=32'd201;
#400 value1=32'd212;value2=32'd230;
#400 value1=32'd233;value2=32'd234;
#400 value1=32'd235;value2=32'd239;
#400 value1=32'd255;value2=32'd257;
#400 value1=32'd297;value2=32'd441;
#400 value1=32'd448;value2=32'd455;
#400 value1=32'd17;value2=32'd63;
#400 value1=32'd202;value2=32'd213;
#400 value1=32'd230;value2=32'd233;
#400 value1=32'd236;value2=32'd237;
#400 value1=32'd240;value2=32'd260;
#400 value1=32'd262;value2=32'd298;
#400 value1=32'd442;value2=32'd449;
#400 value1=32'd64;value2=32'd108;
#400 value1=32'd198;value2=32'd203;
#400 value1=32'd214;value2=32'd231;
#400 value1=32'd232;value2=32'd236;
#400 value1=32'd237;value2=32'd241;
#400 value1=32'd264;value2=32'd266;
#400 value1=32'd299;value2=32'd443;
#400 value1=32'd450;value2=32'd461;
#400 value1=32'd65;value2=32'd204;
#400 value1=32'd209;value2=32'd215;
#400 value1=32'd230;value2=32'd231;
#400 value1=32'd235;value2=32'd236;
#400 value1=32'd242;value2=32'd269;
#400 value1=32'd300;value2=32'd444;
#400 value1=32'd451;value2=32'd462;
#400 value1=32'd66;value2=32'd205;
#400 value1=32'd216;value2=32'd219;
#400 value1=32'd229;value2=32'd230;
#400 value1=32'd231;value2=32'd234;
#400 value1=32'd237;value2=32'd243;
#400 value1=32'd268;value2=32'd271;
#400 value1=32'd301;value2=32'd445;
#400 value1=32'd452;value2=32'd463;
#400 value1=32'd67;value2=32'd206;
#400 value1=32'd209;value2=32'd217;
#400 value1=32'd232;value2=32'd233;
#400 value1=32'd234;value2=32'd237;
#400 value1=32'd244;value2=32'd269;
#400 value1=32'd302;value2=32'd446;
#400 value1=32'd453;value2=32'd464;
#400 value1=32'd68;value2=32'd207;
#400 value1=32'd218;value2=32'd219;
#400 value1=32'd229;value2=32'd232;
#400 value1=32'd233;value2=32'd235;
#400 value1=32'd236;value2=32'd245;
#400 value1=32'd270;value2=32'd273;
#400 value1=32'd303;value2=32'd447;
#400 value1=32'd454;value2=32'd465;
#400 value1=32'd18;value2=32'd69;
#400 value1=32'd200;value2=32'd221;
#400 value1=32'd230;value2=32'd239;
#400 value1=32'd240;value2=32'd242;
#400 value1=32'd243;value2=32'd250;
#400 value1=32'd252;value2=32'd304;
#400 value1=32'd440;value2=32'd477;
#400 value1=32'd70;value2=32'd109;
#400 value1=32'd199;value2=32'd201;
#400 value1=32'd222;value2=32'd231;
#400 value1=32'd238;value2=32'd241;
#400 value1=32'd242;value2=32'd243;
#400 value1=32'd256;value2=32'd258;
#400 value1=32'd305;value2=32'd441;
#400 value1=32'd476;value2=32'd483;
#400 value1=32'd18;value2=32'd71;
#400 value1=32'd202;value2=32'd223;
#400 value1=32'd232;value2=32'd238;
#400 value1=32'd241;value2=32'd244;
#400 value1=32'd245;value2=32'd261;
#400 value1=32'd263;value2=32'd306;
#400 value1=32'd442;value2=32'd477;
#400 value1=32'd72;value2=32'd109;
#400 value1=32'd199;value2=32'd203;
#400 value1=32'd224;value2=32'd233;
#400 value1=32'd239;value2=32'd240;
#400 value1=32'd244;value2=32'd245;
#400 value1=32'd265;value2=32'd267;
#400 value1=32'd307;value2=32'd443;
#400 value1=32'd478;value2=32'd489;
#400 value1=32'd73;value2=32'd204;
#400 value1=32'd210;value2=32'd225;
#400 value1=32'd229;value2=32'd234;
#400 value1=32'd238;value2=32'd239;
#400 value1=32'd243;value2=32'd244;
#400 value1=32'd268;value2=32'd270;
#400 value1=32'd308;value2=32'd444;
#400 value1=32'd479;value2=32'd490;
#400 value1=32'd74;value2=32'd205;
#400 value1=32'd220;value2=32'd226;
#400 value1=32'd235;value2=32'd238;
#400 value1=32'd239;value2=32'd242;
#400 value1=32'd245;value2=32'd272;
#400 value1=32'd309;value2=32'd445;
#400 value1=32'd480;value2=32'd491;
#400 value1=32'd75;value2=32'd206;
#400 value1=32'd210;value2=32'd227;
#400 value1=32'd229;value2=32'd236;
#400 value1=32'd240;value2=32'd241;
#400 value1=32'd242;value2=32'd245;
#400 value1=32'd271;value2=32'd273;
#400 value1=32'd310;value2=32'd446;
#400 value1=32'd481;value2=32'd492;
#400 value1=32'd76;value2=32'd207;
#400 value1=32'd220;value2=32'd228;
#400 value1=32'd237;value2=32'd240;
#400 value1=32'd241;value2=32'd243;
#400 value1=32'd244;value2=32'd272;
#400 value1=32'd311;value2=32'd447;
#400 value1=32'd482;value2=32'd493;
#400 value1=32'd20;value2=32'd77;
#400 value1=32'd110;value2=32'd200;
#400 value1=32'd248;value2=32'd249;
#400 value1=32'd250;value2=32'd253;
#400 value1=32'd255;value2=32'd256;
#400 value1=32'd312;value2=32'd448;
#400 value1=32'd476;value2=32'd504;
#400 value1=32'd19;value2=32'd21;
#400 value1=32'd78;value2=32'd248;
#400 value1=32'd251;value2=32'd252;
#400 value1=32'd253;value2=32'd260;
#400 value1=32'd261;value2=32'd313;
#400 value1=32'd449;value2=32'd477;
#400 value1=32'd22;value2=32'd79;
#400 value1=32'd110;value2=32'd200;
#400 value1=32'd246;value2=32'd247;
#400 value1=32'd251;value2=32'd252;
#400 value1=32'd254;value2=32'd259;
#400 value1=32'd264;value2=32'd265;
#400 value1=32'd314;value2=32'd450;
#400 value1=32'd478;value2=32'd510;
#400 value1=32'd23;value2=32'd80;
#400 value1=32'd211;value2=32'd230;
#400 value1=32'd246;value2=32'd250;
#400 value1=32'd251;value2=32'd255;
#400 value1=32'd260;value2=32'd268;
#400 value1=32'd315;value2=32'd451;
#400 value1=32'd479;value2=32'd511;
#400 value1=32'd24;value2=32'd81;
#400 value1=32'd221;value2=32'd238;
#400 value1=32'd246;value2=32'd249;
#400 value1=32'd252;value2=32'd256;
#400 value1=32'd261;value2=32'd268;
#400 value1=32'd316;value2=32'd452;
#400 value1=32'd480;value2=32'd512;
#400 value1=32'd25;value2=32'd82;
#400 value1=32'd211;value2=32'd230;
#400 value1=32'd247;value2=32'd248;
#400 value1=32'd249;value2=32'd252;
#400 value1=32'd257;value2=32'd262;
#400 value1=32'd269;value2=32'd271;
#400 value1=32'd317;value2=32'd453;
#400 value1=32'd481;value2=32'd513;
#400 value1=32'd26;value2=32'd83;
#400 value1=32'd221;value2=32'd238;
#400 value1=32'd247;value2=32'd248;
#400 value1=32'd250;value2=32'd251;
#400 value1=32'd258;value2=32'd263;
#400 value1=32'd270;value2=32'd272;
#400 value1=32'd318;value2=32'd454;
#400 value1=32'd482;value2=32'd514;
#400 value1=32'd20;value2=32'd84;
#400 value1=32'd112;value2=32'd202;
#400 value1=32'd246;value2=32'd247;
#400 value1=32'd254;value2=32'd257;
#400 value1=32'd258;value2=32'd259;
#400 value1=32'd260;value2=32'd261;
#400 value1=32'd319;value2=32'd455;
#400 value1=32'd483;value2=32'd504;
#400 value1=32'd85;value2=32'd111;
#400 value1=32'd113;value2=32'd201;
#400 value1=32'd203;value2=32'd248;
#400 value1=32'd253;value2=32'd257;
#400 value1=32'd258;value2=32'd264;
#400 value1=32'd265;value2=32'd320;
#400 value1=32'd456;value2=32'd484;
#400 value1=32'd505;value2=32'd525;
#400 value1=32'd86;value2=32'd114;
#400 value1=32'd204;value2=32'd212;
#400 value1=32'd231;value2=32'd246;
#400 value1=32'd249;value2=32'd256;
#400 value1=32'd257;value2=32'd264;
#400 value1=32'd268;value2=32'd321;
#400 value1=32'd457;value2=32'd485;
#400 value1=32'd506;value2=32'd526;
#400 value1=32'd87;value2=32'd115;
#400 value1=32'd205;value2=32'd222;
#400 value1=32'd239;value2=32'd246;
#400 value1=32'd250;value2=32'd255;
#400 value1=32'd258;value2=32'd265;
#400 value1=32'd268;value2=32'd322;
#400 value1=32'd458;value2=32'd486;
#400 value1=32'd507;value2=32'd527;
#400 value1=32'd88;value2=32'd116;
#400 value1=32'd206;value2=32'd212;
#400 value1=32'd231;value2=32'd251;
#400 value1=32'd253;value2=32'd254;
#400 value1=32'd255;value2=32'd258;
#400 value1=32'd266;value2=32'd269;
#400 value1=32'd271;value2=32'd323;
#400 value1=32'd459;value2=32'd487;
#400 value1=32'd508;value2=32'd528;
#400 value1=32'd89;value2=32'd117;
#400 value1=32'd207;value2=32'd222;
#400 value1=32'd239;value2=32'd252;
#400 value1=32'd253;value2=32'd254;
#400 value1=32'd256;value2=32'd257;
#400 value1=32'd267;value2=32'd270;
#400 value1=32'd272;value2=32'd324;
#400 value1=32'd460;value2=32'd488;
#400 value1=32'd509;value2=32'd529;
#400 value1=32'd22;value2=32'd90;
#400 value1=32'd112;value2=32'd202;
#400 value1=32'd248;value2=32'd253;
#400 value1=32'd262;value2=32'd263;
#400 value1=32'd266;value2=32'd267;
#400 value1=32'd325;value2=32'd461;
#400 value1=32'd489;value2=32'd510;
#400 value1=32'd23;value2=32'd91;
#400 value1=32'd213;value2=32'd232;
#400 value1=32'd247;value2=32'd249;
#400 value1=32'd253;value2=32'd261;
#400 value1=32'd262;value2=32'd264;
#400 value1=32'd269;value2=32'd270;
#400 value1=32'd326;value2=32'd462;
#400 value1=32'd490;value2=32'd511;
#400 value1=32'd24;value2=32'd92;
#400 value1=32'd223;value2=32'd240;
#400 value1=32'd247;value2=32'd250;
#400 value1=32'd253;value2=32'd260;
#400 value1=32'd263;value2=32'd265;
#400 value1=32'd271;value2=32'd272;
#400 value1=32'd327;value2=32'd463;
#400 value1=32'd491;value2=32'd512;
#400 value1=32'd25;value2=32'd93;
#400 value1=32'd213;value2=32'd232;
#400 value1=32'd251;value2=32'd259;
#400 value1=32'd260;value2=32'd263;
#400 value1=32'd266;value2=32'd273;
#400 value1=32'd328;value2=32'd464;
#400 value1=32'd492;value2=32'd513;
#400 value1=32'd26;value2=32'd94;
#400 value1=32'd223;value2=32'd240;
#400 value1=32'd252;value2=32'd259;
#400 value1=32'd261;value2=32'd262;
#400 value1=32'd267;value2=32'd273;
#400 value1=32'd329;value2=32'd465;
#400 value1=32'd493;value2=32'd514;
#400 value1=32'd95;value2=32'd114;
#400 value1=32'd204;value2=32'd214;
#400 value1=32'd233;value2=32'd248;
#400 value1=32'd254;value2=32'd255;
#400 value1=32'd260;value2=32'd265;
#400 value1=32'd266;value2=32'd269;
#400 value1=32'd270;value2=32'd330;
#400 value1=32'd466;value2=32'd494;
#400 value1=32'd515;value2=32'd540;
#400 value1=32'd96;value2=32'd115;
#400 value1=32'd205;value2=32'd224;
#400 value1=32'd241;value2=32'd248;
#400 value1=32'd254;value2=32'd256;
#400 value1=32'd261;value2=32'd264;
#400 value1=32'd267;value2=32'd271;
#400 value1=32'd272;value2=32'd331;
#400 value1=32'd467;value2=32'd495;
#400 value1=32'd516;value2=32'd541;
#400 value1=32'd97;value2=32'd116;
#400 value1=32'd206;value2=32'd214;
#400 value1=32'd233;value2=32'd257;
#400 value1=32'd259;value2=32'd262;
#400 value1=32'd264;value2=32'd267;
#400 value1=32'd273;value2=32'd332;
#400 value1=32'd468;value2=32'd496;
#400 value1=32'd517;value2=32'd542;
#400 value1=32'd98;value2=32'd117;
#400 value1=32'd207;value2=32'd224;
#400 value1=32'd241;value2=32'd258;
#400 value1=32'd259;value2=32'd263;
#400 value1=32'd265;value2=32'd266;
#400 value1=32'd273;value2=32'd333;
#400 value1=32'd469;value2=32'd497;
#400 value1=32'd518;value2=32'd543;
#400 value1=32'd99;value2=32'd216;
#400 value1=32'd225;value2=32'd235;
#400 value1=32'd242;value2=32'd249;
#400 value1=32'd250;value2=32'd255;
#400 value1=32'd256;value2=32'd270;
#400 value1=32'd271;value2=32'd334;
#400 value1=32'd470;value2=32'd498;
#400 value1=32'd519;value2=32'd544;
#400 value1=32'd100;value2=32'd215;
#400 value1=32'd217;value2=32'd234;
#400 value1=32'd236;value2=32'd251;
#400 value1=32'd257;value2=32'd260;
#400 value1=32'd264;value2=32'd270;
#400 value1=32'd271;value2=32'd335;
#400 value1=32'd471;value2=32'd499;
#400 value1=32'd520;value2=32'd545;
#400 value1=32'd101;value2=32'd218;
#400 value1=32'd225;value2=32'd237;
#400 value1=32'd242;value2=32'd252;
#400 value1=32'd258;value2=32'd260;
#400 value1=32'd264;value2=32'd268;
#400 value1=32'd269;value2=32'd272;
#400 value1=32'd273;value2=32'd336;
#400 value1=32'd472;value2=32'd500;
#400 value1=32'd521;value2=32'd546;
#400 value1=32'd102;value2=32'd216;
#400 value1=32'd227;value2=32'd235;
#400 value1=32'd244;value2=32'd251;
#400 value1=32'd257;value2=32'd261;
#400 value1=32'd265;value2=32'd268;
#400 value1=32'd269;value2=32'd272;
#400 value1=32'd273;value2=32'd337;
#400 value1=32'd473;value2=32'd501;
#400 value1=32'd522;value2=32'd547;
#400 value1=32'd103;value2=32'd226;
#400 value1=32'd228;value2=32'd243;
#400 value1=32'd245;value2=32'd252;
#400 value1=32'd258;value2=32'd261;
#400 value1=32'd265;value2=32'd270;
#400 value1=32'd271;value2=32'd338;
#400 value1=32'd474;value2=32'd502;
#400 value1=32'd523;value2=32'd548;
#400 value1=32'd104;value2=32'd218;
#400 value1=32'd227;value2=32'd237;
#400 value1=32'd244;value2=32'd262;
#400 value1=32'd263;value2=32'd266;
#400 value1=32'd267;value2=32'd270;
#400 value1=32'd271;value2=32'd339;
#400 value1=32'd475;value2=32'd503;
#400 value1=32'd524;value2=32'd549;
#400 value1=32'd27;value2=32'd28;
#400 value1=32'd118;value2=32'd119;
#400 value1=32'd130;value2=32'd208;
#400 value1=32'd276;value2=32'd282;
#400 value1=32'd284;value2=32'd285;
#400 value1=32'd291;value2=32'd293;
#400 value1=32'd340;value2=32'd341;
#400 value1=32'd343;value2=32'd345;
#400 value1=32'd29;value2=32'd120;
#400 value1=32'd131;value2=32'd196;
#400 value1=32'd209;value2=32'd276;
#400 value1=32'd281;value2=32'd283;
#400 value1=32'd285;value2=32'd300;
#400 value1=32'd302;value2=32'd350;
#400 value1=32'd352;value2=32'd354;
#400 value1=32'd30;value2=32'd121;
#400 value1=32'd132;value2=32'd196;
#400 value1=32'd210;value2=32'd274;
#400 value1=32'd275;value2=32'd282;
#400 value1=32'd284;value2=32'd286;
#400 value1=32'd295;value2=32'd308;
#400 value1=32'd310;value2=32'd350;
#400 value1=32'd360;value2=32'd362;
#400 value1=32'd27;value2=32'd31;
#400 value1=32'd122;value2=32'd133;
#400 value1=32'd196;value2=32'd211;
#400 value1=32'd278;value2=32'd279;
#400 value1=32'd281;value2=32'd282;
#400 value1=32'd287;value2=32'd296;
#400 value1=32'd315;value2=32'd317;
#400 value1=32'd351;value2=32'd359;
#400 value1=32'd367;value2=32'd369;
#400 value1=32'd32;value2=32'd118;
#400 value1=32'd123;value2=32'd134;
#400 value1=32'd212;value2=32'd277;
#400 value1=32'd280;value2=32'd281;
#400 value1=32'd282;value2=32'd288;
#400 value1=32'd297;value2=32'd321;
#400 value1=32'd323;value2=32'd352;
#400 value1=32'd360;value2=32'd375;
#400 value1=32'd27;value2=32'd33;
#400 value1=32'd124;value2=32'd135;
#400 value1=32'd196;value2=32'd213;
#400 value1=32'd277;value2=32'd280;
#400 value1=32'd283;value2=32'd284;
#400 value1=32'd289;value2=32'd298;
#400 value1=32'd326;value2=32'd328;
#400 value1=32'd353;value2=32'd361;
#400 value1=32'd374;value2=32'd380;
#400 value1=32'd34;value2=32'd118;
#400 value1=32'd125;value2=32'd136;
#400 value1=32'd214;value2=32'd278;
#400 value1=32'd279;value2=32'd283;
#400 value1=32'd284;value2=32'd290;
#400 value1=32'd299;value2=32'd330;
#400 value1=32'd332;value2=32'd354;
#400 value1=32'd362;value2=32'd375;
#400 value1=32'd35;value2=32'd126;
#400 value1=32'd137;value2=32'd215;
#400 value1=32'd275;value2=32'd277;
#400 value1=32'd278;value2=32'd282;
#400 value1=32'd283;value2=32'd291;
#400 value1=32'd300;value2=32'd335;
#400 value1=32'd355;value2=32'd363;
#400 value1=32'd376;value2=32'd385;
#400 value1=32'd36;value2=32'd127;
#400 value1=32'd138;value2=32'd216;
#400 value1=32'd274;value2=32'd276;
#400 value1=32'd277;value2=32'd278;
#400 value1=32'd281;value2=32'd284;
#400 value1=32'd292;value2=32'd301;
#400 value1=32'd334;value2=32'd337;
#400 value1=32'd356;value2=32'd364;
#400 value1=32'd377;value2=32'd386;
#400 value1=32'd37;value2=32'd128;
#400 value1=32'd139;value2=32'd217;
#400 value1=32'd275;value2=32'd279;
#400 value1=32'd280;value2=32'd281;
#400 value1=32'd284;value2=32'd293;
#400 value1=32'd302;value2=32'd335;
#400 value1=32'd357;value2=32'd365;
#400 value1=32'd378;value2=32'd387;
#400 value1=32'd38;value2=32'd129;
#400 value1=32'd140;value2=32'd218;
#400 value1=32'd274;value2=32'd276;
#400 value1=32'd279;value2=32'd280;
#400 value1=32'd282;value2=32'd283;
#400 value1=32'd294;value2=32'd303;
#400 value1=32'd336;value2=32'd339;
#400 value1=32'd358;value2=32'd366;
#400 value1=32'd379;value2=32'd388;
#400 value1=32'd29;value2=32'd120;
#400 value1=32'd141;value2=32'd197;
#400 value1=32'd219;value2=32'd274;
#400 value1=32'd275;value2=32'd286;
#400 value1=32'd291;value2=32'd293;
#400 value1=32'd295;value2=32'd301;
#400 value1=32'd303;value2=32'd395;
#400 value1=32'd397;value2=32'd399;
#400 value1=32'd30;value2=32'd121;
#400 value1=32'd142;value2=32'd197;
#400 value1=32'd220;value2=32'd276;
#400 value1=32'd285;value2=32'd292;
#400 value1=32'd294;value2=32'd309;
#400 value1=32'd311;value2=32'd395;
#400 value1=32'd405;value2=32'd407;
#400 value1=32'd28;value2=32'd31;
#400 value1=32'd122;value2=32'd143;
#400 value1=32'd197;value2=32'd221;
#400 value1=32'd277;value2=32'd288;
#400 value1=32'd289;value2=32'd291;
#400 value1=32'd292;value2=32'd304;
#400 value1=32'd316;value2=32'd318;
#400 value1=32'd396;value2=32'd404;
#400 value1=32'd412;value2=32'd414;
#400 value1=32'd32;value2=32'd119;
#400 value1=32'd123;value2=32'd144;
#400 value1=32'd222;value2=32'd278;
#400 value1=32'd287;value2=32'd290;
#400 value1=32'd291;value2=32'd292;
#400 value1=32'd305;value2=32'd322;
#400 value1=32'd324;value2=32'd397;
#400 value1=32'd405;value2=32'd420;
#400 value1=32'd28;value2=32'd33;
#400 value1=32'd124;value2=32'd145;
#400 value1=32'd197;value2=32'd223;
#400 value1=32'd279;value2=32'd287;
#400 value1=32'd290;value2=32'd293;
#400 value1=32'd294;value2=32'd306;
#400 value1=32'd327;value2=32'd329;
#400 value1=32'd398;value2=32'd406;
#400 value1=32'd419;value2=32'd425;
#400 value1=32'd34;value2=32'd119;
#400 value1=32'd125;value2=32'd146;
#400 value1=32'd224;value2=32'd280;
#400 value1=32'd288;value2=32'd289;
#400 value1=32'd293;value2=32'd294;
#400 value1=32'd307;value2=32'd331;
#400 value1=32'd333;value2=32'd399;
#400 value1=32'd407;value2=32'd420;
#400 value1=32'd35;value2=32'd126;
#400 value1=32'd147;value2=32'd225;
#400 value1=32'd274;value2=32'd281;
#400 value1=32'd285;value2=32'd287;
#400 value1=32'd288;value2=32'd292;
#400 value1=32'd293;value2=32'd308;
#400 value1=32'd334;value2=32'd336;
#400 value1=32'd400;value2=32'd408;
#400 value1=32'd421;value2=32'd430;
#400 value1=32'd36;value2=32'd127;
#400 value1=32'd148;value2=32'd226;
#400 value1=32'd282;value2=32'd286;
#400 value1=32'd287;value2=32'd288;
#400 value1=32'd291;value2=32'd294;
#400 value1=32'd309;value2=32'd338;
#400 value1=32'd401;value2=32'd409;
#400 value1=32'd422;value2=32'd431;
#400 value1=32'd37;value2=32'd128;
#400 value1=32'd149;value2=32'd227;
#400 value1=32'd274;value2=32'd283;
#400 value1=32'd285;value2=32'd289;
#400 value1=32'd290;value2=32'd291;
#400 value1=32'd294;value2=32'd310;
#400 value1=32'd337;value2=32'd339;
#400 value1=32'd402;value2=32'd410;
#400 value1=32'd423;value2=32'd432;
#400 value1=32'd38;value2=32'd129;
#400 value1=32'd150;value2=32'd228;
#400 value1=32'd284;value2=32'd286;
#400 value1=32'd289;value2=32'd290;
#400 value1=32'd292;value2=32'd293;
#400 value1=32'd311;value2=32'd338;
#400 value1=32'd403;value2=32'd411;
#400 value1=32'd424;value2=32'd433;
#400 value1=32'd151;value2=32'd198;
#400 value1=32'd199;value2=32'd229;
#400 value1=32'd276;value2=32'd285;
#400 value1=32'd301;value2=32'd303;
#400 value1=32'd308;value2=32'd310;
#400 value1=32'd441;value2=32'd443;
#400 value1=32'd29;value2=32'd152;
#400 value1=32'd198;value2=32'd200;
#400 value1=32'd230;value2=32'd277;
#400 value1=32'd297;value2=32'd298;
#400 value1=32'd300;value2=32'd301;
#400 value1=32'd304;value2=32'd315;
#400 value1=32'd317;value2=32'd440;
#400 value1=32'd448;value2=32'd450;
#400 value1=32'd120;value2=32'd153;
#400 value1=32'd201;value2=32'd231;
#400 value1=32'd278;value2=32'd296;
#400 value1=32'd299;value2=32'd300;
#400 value1=32'd301;value2=32'd305;
#400 value1=32'd321;value2=32'd323;
#400 value1=32'd441;value2=32'd456;
#400 value1=32'd29;value2=32'd154;
#400 value1=32'd198;value2=32'd202;
#400 value1=32'd232;value2=32'd279;
#400 value1=32'd296;value2=32'd299;
#400 value1=32'd302;value2=32'd303;
#400 value1=32'd306;value2=32'd326;
#400 value1=32'd328;value2=32'd442;
#400 value1=32'd455;value2=32'd461;
#400 value1=32'd120;value2=32'd155;
#400 value1=32'd203;value2=32'd233;
#400 value1=32'd280;value2=32'd297;
#400 value1=32'd298;value2=32'd302;
#400 value1=32'd303;value2=32'd307;
#400 value1=32'd330;value2=32'd332;
#400 value1=32'd443;value2=32'd456;
#400 value1=32'd156;value2=32'd204;
#400 value1=32'd234;value2=32'd275;
#400 value1=32'd281;value2=32'd296;
#400 value1=32'd297;value2=32'd301;
#400 value1=32'd302;value2=32'd308;
#400 value1=32'd335;value2=32'd444;
#400 value1=32'd457;value2=32'd466;
#400 value1=32'd157;value2=32'd205;
#400 value1=32'd235;value2=32'd282;
#400 value1=32'd285;value2=32'd295;
#400 value1=32'd296;value2=32'd297;
#400 value1=32'd300;value2=32'd303;
#400 value1=32'd309;value2=32'd334;
#400 value1=32'd337;value2=32'd445;
#400 value1=32'd458;value2=32'd467;
#400 value1=32'd158;value2=32'd206;
#400 value1=32'd236;value2=32'd275;
#400 value1=32'd283;value2=32'd298;
#400 value1=32'd299;value2=32'd300;
#400 value1=32'd303;value2=32'd310;
#400 value1=32'd335;value2=32'd446;
#400 value1=32'd459;value2=32'd468;
#400 value1=32'd159;value2=32'd207;
#400 value1=32'd237;value2=32'd284;
#400 value1=32'd285;value2=32'd295;
#400 value1=32'd298;value2=32'd299;
#400 value1=32'd301;value2=32'd302;
#400 value1=32'd311;value2=32'd336;
#400 value1=32'd339;value2=32'd447;
#400 value1=32'd460;value2=32'd469;
#400 value1=32'd30;value2=32'd160;
#400 value1=32'd199;value2=32'd200;
#400 value1=32'd238;value2=32'd287;
#400 value1=32'd296;value2=32'd305;
#400 value1=32'd306;value2=32'd308;
#400 value1=32'd309;value2=32'd316;
#400 value1=32'd318;value2=32'd440;
#400 value1=32'd476;value2=32'd478;
#400 value1=32'd121;value2=32'd161;
#400 value1=32'd201;value2=32'd239;
#400 value1=32'd288;value2=32'd297;
#400 value1=32'd304;value2=32'd307;
#400 value1=32'd308;value2=32'd309;
#400 value1=32'd322;value2=32'd324;
#400 value1=32'd441;value2=32'd484;
#400 value1=32'd30;value2=32'd162;
#400 value1=32'd199;value2=32'd202;
#400 value1=32'd240;value2=32'd289;
#400 value1=32'd298;value2=32'd304;
#400 value1=32'd307;value2=32'd310;
#400 value1=32'd311;value2=32'd327;
#400 value1=32'd329;value2=32'd442;
#400 value1=32'd483;value2=32'd489;
#400 value1=32'd121;value2=32'd163;
#400 value1=32'd203;value2=32'd241;
#400 value1=32'd290;value2=32'd299;
#400 value1=32'd305;value2=32'd306;
#400 value1=32'd310;value2=32'd311;
#400 value1=32'd331;value2=32'd333;
#400 value1=32'd443;value2=32'd484;
#400 value1=32'd164;value2=32'd204;
#400 value1=32'd242;value2=32'd276;
#400 value1=32'd291;value2=32'd295;
#400 value1=32'd300;value2=32'd304;
#400 value1=32'd305;value2=32'd309;
#400 value1=32'd310;value2=32'd334;
#400 value1=32'd336;value2=32'd444;
#400 value1=32'd485;value2=32'd494;
#400 value1=32'd165;value2=32'd205;
#400 value1=32'd243;value2=32'd286;
#400 value1=32'd292;value2=32'd301;
#400 value1=32'd304;value2=32'd305;
#400 value1=32'd308;value2=32'd311;
#400 value1=32'd338;value2=32'd445;
#400 value1=32'd486;value2=32'd495;
#400 value1=32'd166;value2=32'd206;
#400 value1=32'd244;value2=32'd276;
#400 value1=32'd293;value2=32'd295;
#400 value1=32'd302;value2=32'd306;
#400 value1=32'd307;value2=32'd308;
#400 value1=32'd311;value2=32'd337;
#400 value1=32'd339;value2=32'd446;
#400 value1=32'd487;value2=32'd496;
#400 value1=32'd167;value2=32'd207;
#400 value1=32'd245;value2=32'd286;
#400 value1=32'd294;value2=32'd303;
#400 value1=32'd306;value2=32'd307;
#400 value1=32'd309;value2=32'd310;
#400 value1=32'd338;value2=32'd447;
#400 value1=32'd488;value2=32'd497;
#400 value1=32'd32;value2=32'd122;
#400 value1=32'd168;value2=32'd201;
#400 value1=32'd246;value2=32'd314;
#400 value1=32'd315;value2=32'd316;
#400 value1=32'd319;value2=32'd321;
#400 value1=32'd322;value2=32'd448;
#400 value1=32'd476;value2=32'd505;
#400 value1=32'd31;value2=32'd33;
#400 value1=32'd169;value2=32'd200;
#400 value1=32'd202;value2=32'd247;
#400 value1=32'd314;value2=32'd317;
#400 value1=32'd318;value2=32'd319;
#400 value1=32'd326;value2=32'd327;
#400 value1=32'd449;value2=32'd477;
#400 value1=32'd504;value2=32'd510;
#400 value1=32'd34;value2=32'd122;
#400 value1=32'd170;value2=32'd203;
#400 value1=32'd248;value2=32'd312;
#400 value1=32'd313;value2=32'd317;
#400 value1=32'd318;value2=32'd320;
#400 value1=32'd325;value2=32'd330;
#400 value1=32'd331;value2=32'd450;
#400 value1=32'd478;value2=32'd505;
#400 value1=32'd35;value2=32'd171;
#400 value1=32'd204;value2=32'd249;
#400 value1=32'd277;value2=32'd296;
#400 value1=32'd312;value2=32'd316;
#400 value1=32'd317;value2=32'd321;
#400 value1=32'd326;value2=32'd334;
#400 value1=32'd451;value2=32'd479;
#400 value1=32'd506;value2=32'd515;
#400 value1=32'd36;value2=32'd172;
#400 value1=32'd205;value2=32'd250;
#400 value1=32'd287;value2=32'd304;
#400 value1=32'd312;value2=32'd315;
#400 value1=32'd318;value2=32'd322;
#400 value1=32'd327;value2=32'd334;
#400 value1=32'd452;value2=32'd480;
#400 value1=32'd507;value2=32'd516;
#400 value1=32'd37;value2=32'd173;
#400 value1=32'd206;value2=32'd251;
#400 value1=32'd277;value2=32'd296;
#400 value1=32'd313;value2=32'd314;
#400 value1=32'd315;value2=32'd318;
#400 value1=32'd323;value2=32'd328;
#400 value1=32'd335;value2=32'd337;
#400 value1=32'd453;value2=32'd481;
#400 value1=32'd508;value2=32'd517;
#400 value1=32'd38;value2=32'd174;
#400 value1=32'd207;value2=32'd252;
#400 value1=32'd287;value2=32'd304;
#400 value1=32'd313;value2=32'd314;
#400 value1=32'd316;value2=32'd317;
#400 value1=32'd324;value2=32'd329;
#400 value1=32'd336;value2=32'd338;
#400 value1=32'd454;value2=32'd482;
#400 value1=32'd509;value2=32'd518;
#400 value1=32'd32;value2=32'd124;
#400 value1=32'd175;value2=32'd201;
#400 value1=32'd253;value2=32'd312;
#400 value1=32'd313;value2=32'd320;
#400 value1=32'd323;value2=32'd324;
#400 value1=32'd325;value2=32'd326;
#400 value1=32'd327;value2=32'd455;
#400 value1=32'd483;value2=32'd525;
#400 value1=32'd123;value2=32'd125;
#400 value1=32'd176;value2=32'd254;
#400 value1=32'd314;value2=32'd319;
#400 value1=32'd323;value2=32'd324;
#400 value1=32'd330;value2=32'd331;
#400 value1=32'd456;value2=32'd484;
#400 value1=32'd126;value2=32'd177;
#400 value1=32'd255;value2=32'd278;
#400 value1=32'd297;value2=32'd312;
#400 value1=32'd315;value2=32'd322;
#400 value1=32'd323;value2=32'd330;
#400 value1=32'd334;value2=32'd457;
#400 value1=32'd485;value2=32'd530;
#400 value1=32'd127;value2=32'd178;
#400 value1=32'd256;value2=32'd288;
#400 value1=32'd305;value2=32'd312;
#400 value1=32'd316;value2=32'd321;
#400 value1=32'd324;value2=32'd331;
#400 value1=32'd334;value2=32'd458;
#400 value1=32'd486;value2=32'd531;
#400 value1=32'd128;value2=32'd179;
#400 value1=32'd257;value2=32'd278;
#400 value1=32'd297;value2=32'd317;
#400 value1=32'd319;value2=32'd320;
#400 value1=32'd321;value2=32'd324;
#400 value1=32'd332;value2=32'd335;
#400 value1=32'd337;value2=32'd459;
#400 value1=32'd487;value2=32'd532;
#400 value1=32'd129;value2=32'd180;
#400 value1=32'd258;value2=32'd288;
#400 value1=32'd305;value2=32'd318;
#400 value1=32'd319;value2=32'd320;
#400 value1=32'd322;value2=32'd323;
#400 value1=32'd333;value2=32'd336;
#400 value1=32'd338;value2=32'd460;
#400 value1=32'd488;value2=32'd533;
#400 value1=32'd34;value2=32'd124;
#400 value1=32'd181;value2=32'd203;
#400 value1=32'd259;value2=32'd314;
#400 value1=32'd319;value2=32'd328;
#400 value1=32'd329;value2=32'd332;
#400 value1=32'd333;value2=32'd461;
#400 value1=32'd489;value2=32'd525;
#400 value1=32'd35;value2=32'd182;
#400 value1=32'd204;value2=32'd260;
#400 value1=32'd279;value2=32'd298;
#400 value1=32'd313;value2=32'd315;
#400 value1=32'd319;value2=32'd327;
#400 value1=32'd328;value2=32'd330;
#400 value1=32'd335;value2=32'd336;
#400 value1=32'd462;value2=32'd490;
#400 value1=32'd526;value2=32'd540;
#400 value1=32'd36;value2=32'd183;
#400 value1=32'd205;value2=32'd261;
#400 value1=32'd289;value2=32'd306;
#400 value1=32'd313;value2=32'd316;
#400 value1=32'd319;value2=32'd326;
#400 value1=32'd329;value2=32'd331;
#400 value1=32'd337;value2=32'd338;
#400 value1=32'd463;value2=32'd491;
#400 value1=32'd527;value2=32'd541;
#400 value1=32'd37;value2=32'd184;
#400 value1=32'd206;value2=32'd262;
#400 value1=32'd279;value2=32'd298;
#400 value1=32'd317;value2=32'd325;
#400 value1=32'd326;value2=32'd329;
#400 value1=32'd332;value2=32'd339;
#400 value1=32'd464;value2=32'd492;
#400 value1=32'd528;value2=32'd542;
#400 value1=32'd38;value2=32'd185;
#400 value1=32'd207;value2=32'd263;
#400 value1=32'd289;value2=32'd306;
#400 value1=32'd318;value2=32'd325;
#400 value1=32'd327;value2=32'd328;
#400 value1=32'd333;value2=32'd339;
#400 value1=32'd465;value2=32'd493;
#400 value1=32'd529;value2=32'd543;
#400 value1=32'd126;value2=32'd186;
#400 value1=32'd264;value2=32'd280;
#400 value1=32'd299;value2=32'd314;
#400 value1=32'd320;value2=32'd321;
#400 value1=32'd326;value2=32'd331;
#400 value1=32'd332;value2=32'd335;
#400 value1=32'd336;value2=32'd466;
#400 value1=32'd494;value2=32'd530;
#400 value1=32'd127;value2=32'd187;
#400 value1=32'd265;value2=32'd290;
#400 value1=32'd307;value2=32'd314;
#400 value1=32'd320;value2=32'd322;
#400 value1=32'd327;value2=32'd330;
#400 value1=32'd333;value2=32'd337;
#400 value1=32'd338;value2=32'd467;
#400 value1=32'd495;value2=32'd531;
#400 value1=32'd128;value2=32'd188;
#400 value1=32'd266;value2=32'd280;
#400 value1=32'd299;value2=32'd323;
#400 value1=32'd325;value2=32'd328;
#400 value1=32'd330;value2=32'd333;
#400 value1=32'd339;value2=32'd468;
#400 value1=32'd496;value2=32'd532;
#400 value1=32'd129;value2=32'd189;
#400 value1=32'd267;value2=32'd290;
#400 value1=32'd307;value2=32'd324;
#400 value1=32'd325;value2=32'd329;
#400 value1=32'd331;value2=32'd332;
#400 value1=32'd339;value2=32'd469;
#400 value1=32'd497;value2=32'd533;
#400 value1=32'd190;value2=32'd268;
#400 value1=32'd282;value2=32'd291;
#400 value1=32'd301;value2=32'd308;
#400 value1=32'd315;value2=32'd316;
#400 value1=32'd321;value2=32'd322;
#400 value1=32'd336;value2=32'd337;
#400 value1=32'd470;value2=32'd498;
#400 value1=32'd534;value2=32'd550;
#400 value1=32'd191;value2=32'd269;
#400 value1=32'd281;value2=32'd283;
#400 value1=32'd300;value2=32'd302;
#400 value1=32'd317;value2=32'd323;
#400 value1=32'd326;value2=32'd330;
#400 value1=32'd336;value2=32'd337;
#400 value1=32'd471;value2=32'd499;
#400 value1=32'd535;value2=32'd551;
#400 value1=32'd192;value2=32'd270;
#400 value1=32'd284;value2=32'd291;
#400 value1=32'd303;value2=32'd308;
#400 value1=32'd318;value2=32'd324;
#400 value1=32'd326;value2=32'd330;
#400 value1=32'd334;value2=32'd335;
#400 value1=32'd338;value2=32'd339;
#400 value1=32'd472;value2=32'd500;
#400 value1=32'd536;value2=32'd552;
#400 value1=32'd193;value2=32'd271;
#400 value1=32'd282;value2=32'd293;
#400 value1=32'd301;value2=32'd310;
#400 value1=32'd317;value2=32'd323;
#400 value1=32'd327;value2=32'd331;
#400 value1=32'd334;value2=32'd335;
#400 value1=32'd338;value2=32'd339;
#400 value1=32'd473;value2=32'd501;
#400 value1=32'd537;value2=32'd553;
#400 value1=32'd194;value2=32'd272;
#400 value1=32'd292;value2=32'd294;
#400 value1=32'd309;value2=32'd311;
#400 value1=32'd318;value2=32'd324;
#400 value1=32'd327;value2=32'd331;
#400 value1=32'd336;value2=32'd337;
#400 value1=32'd474;value2=32'd502;
#400 value1=32'd538;value2=32'd554;
#400 value1=32'd195;value2=32'd273;
#400 value1=32'd284;value2=32'd293;
#400 value1=32'd303;value2=32'd310;
#400 value1=32'd328;value2=32'd329;
#400 value1=32'd332;value2=32'd333;
#400 value1=32'd336;value2=32'd337;
#400 value1=32'd475;value2=32'd503;
#400 value1=32'd539;value2=32'd555;
#400 value1=32'd40;value2=32'd50;
#400 value1=32'd131;value2=32'd141;
#400 value1=32'd208;value2=32'd274;
#400 value1=32'd341;value2=32'd346;
#400 value1=32'd348;value2=32'd350;
#400 value1=32'd356;value2=32'd358;
#400 value1=32'd400;value2=32'd402;
#400 value1=32'd41;value2=32'd51;
#400 value1=32'd132;value2=32'd142;
#400 value1=32'd208;value2=32'd274;
#400 value1=32'd340;value2=32'd347;
#400 value1=32'd349;value2=32'd364;
#400 value1=32'd366;value2=32'd395;
#400 value1=32'd408;value2=32'd410;
#400 value1=32'd39;value2=32'd42;
#400 value1=32'd52;value2=32'd133;
#400 value1=32'd143;value2=32'd208;
#400 value1=32'd343;value2=32'd344;
#400 value1=32'd346;value2=32'd347;
#400 value1=32'd359;value2=32'd371;
#400 value1=32'd373;value2=32'd396;
#400 value1=32'd415;value2=32'd417;
#400 value1=32'd43;value2=32'd53;
#400 value1=32'd130;value2=32'd134;
#400 value1=32'd144;value2=32'd274;
#400 value1=32'd342;value2=32'd345;
#400 value1=32'd346;value2=32'd347;
#400 value1=32'd360;value2=32'd377;
#400 value1=32'd379;value2=32'd397;
#400 value1=32'd421;value2=32'd423;
#400 value1=32'd39;value2=32'd44;
#400 value1=32'd54;value2=32'd135;
#400 value1=32'd145;value2=32'd208;
#400 value1=32'd342;value2=32'd345;
#400 value1=32'd348;value2=32'd349;
#400 value1=32'd361;value2=32'd382;
#400 value1=32'd384;value2=32'd398;
#400 value1=32'd426;value2=32'd428;
#400 value1=32'd45;value2=32'd55;
#400 value1=32'd130;value2=32'd136;
#400 value1=32'd146;value2=32'd274;
#400 value1=32'd343;value2=32'd344;
#400 value1=32'd348;value2=32'd349;
#400 value1=32'd362;value2=32'd386;
#400 value1=32'd388;value2=32'd399;
#400 value1=32'd430;value2=32'd432;
#400 value1=32'd46;value2=32'd56;
#400 value1=32'd137;value2=32'd147;
#400 value1=32'd340;value2=32'd342;
#400 value1=32'd343;value2=32'd347;
#400 value1=32'd348;value2=32'd363;
#400 value1=32'd389;value2=32'd391;
#400 value1=32'd400;value2=32'd435;
#400 value1=32'd47;value2=32'd57;
#400 value1=32'd138;value2=32'd148;
#400 value1=32'd341;value2=32'd342;
#400 value1=32'd343;value2=32'd346;
#400 value1=32'd349;value2=32'd364;
#400 value1=32'd393;value2=32'd401;
#400 value1=32'd434;value2=32'd437;
#400 value1=32'd48;value2=32'd58;
#400 value1=32'd139;value2=32'd149;
#400 value1=32'd340;value2=32'd344;
#400 value1=32'd345;value2=32'd346;
#400 value1=32'd349;value2=32'd365;
#400 value1=32'd392;value2=32'd394;
#400 value1=32'd402;value2=32'd435;
#400 value1=32'd49;value2=32'd59;
#400 value1=32'd140;value2=32'd150;
#400 value1=32'd341;value2=32'd344;
#400 value1=32'd345;value2=32'd347;
#400 value1=32'd348;value2=32'd366;
#400 value1=32'd393;value2=32'd403;
#400 value1=32'd436;value2=32'd439;
#400 value1=32'd60;value2=32'd151;
#400 value1=32'd209;value2=32'd210;
#400 value1=32'd275;value2=32'd276;
#400 value1=32'd340;value2=32'd356;
#400 value1=32'd358;value2=32'd363;
#400 value1=32'd365;value2=32'd395;
#400 value1=32'd444;value2=32'd446;
#400 value1=32'd40;value2=32'd61;
#400 value1=32'd152;value2=32'd209;
#400 value1=32'd211;value2=32'd277;
#400 value1=32'd352;value2=32'd353;
#400 value1=32'd355;value2=32'd356;
#400 value1=32'd359;value2=32'd370;
#400 value1=32'd372;value2=32'd396;
#400 value1=32'd451;value2=32'd453;
#400 value1=32'd62;value2=32'd131;
#400 value1=32'd153;value2=32'd212;
#400 value1=32'd275;value2=32'd278;
#400 value1=32'd351;value2=32'd354;
#400 value1=32'd355;value2=32'd356;
#400 value1=32'd360;value2=32'd376;
#400 value1=32'd378;value2=32'd397;
#400 value1=32'd457;value2=32'd459;
#400 value1=32'd40;value2=32'd63;
#400 value1=32'd154;value2=32'd209;
#400 value1=32'd213;value2=32'd279;
#400 value1=32'd351;value2=32'd354;
#400 value1=32'd357;value2=32'd358;
#400 value1=32'd361;value2=32'd381;
#400 value1=32'd383;value2=32'd398;
#400 value1=32'd462;value2=32'd464;
#400 value1=32'd64;value2=32'd131;
#400 value1=32'd155;value2=32'd214;
#400 value1=32'd275;value2=32'd280;
#400 value1=32'd352;value2=32'd353;
#400 value1=32'd357;value2=32'd358;
#400 value1=32'd362;value2=32'd385;
#400 value1=32'd387;value2=32'd399;
#400 value1=32'd466;value2=32'd468;
#400 value1=32'd65;value2=32'd156;
#400 value1=32'd215;value2=32'd281;
#400 value1=32'd351;value2=32'd352;
#400 value1=32'd356;value2=32'd357;
#400 value1=32'd363;value2=32'd390;
#400 value1=32'd400;value2=32'd471;
#400 value1=32'd66;value2=32'd157;
#400 value1=32'd216;value2=32'd282;
#400 value1=32'd340;value2=32'd350;
#400 value1=32'd351;value2=32'd352;
#400 value1=32'd355;value2=32'd358;
#400 value1=32'd364;value2=32'd389;
#400 value1=32'd392;value2=32'd401;
#400 value1=32'd470;value2=32'd473;
#400 value1=32'd67;value2=32'd158;
#400 value1=32'd217;value2=32'd283;
#400 value1=32'd353;value2=32'd354;
#400 value1=32'd355;value2=32'd358;
#400 value1=32'd365;value2=32'd390;
#400 value1=32'd402;value2=32'd471;
#400 value1=32'd68;value2=32'd159;
#400 value1=32'd218;value2=32'd284;
#400 value1=32'd340;value2=32'd350;
#400 value1=32'd353;value2=32'd354;
#400 value1=32'd356;value2=32'd357;
#400 value1=32'd366;value2=32'd391;
#400 value1=32'd394;value2=32'd403;
#400 value1=32'd472;value2=32'd475;
#400 value1=32'd41;value2=32'd69;
#400 value1=32'd160;value2=32'd210;
#400 value1=32'd211;value2=32'd277;
#400 value1=32'd342;value2=32'd351;
#400 value1=32'd360;value2=32'd361;
#400 value1=32'd363;value2=32'd364;
#400 value1=32'd371;value2=32'd373;
#400 value1=32'd404;value2=32'd440;
#400 value1=32'd479;value2=32'd481;
#400 value1=32'd70;value2=32'd132;
#400 value1=32'd161;value2=32'd212;
#400 value1=32'd276;value2=32'd278;
#400 value1=32'd343;value2=32'd352;
#400 value1=32'd359;value2=32'd362;
#400 value1=32'd363;value2=32'd364;
#400 value1=32'd377;value2=32'd379;
#400 value1=32'd405;value2=32'd441;
#400 value1=32'd485;value2=32'd487;
#400 value1=32'd41;value2=32'd71;
#400 value1=32'd162;value2=32'd210;
#400 value1=32'd213;value2=32'd279;
#400 value1=32'd344;value2=32'd353;
#400 value1=32'd359;value2=32'd362;
#400 value1=32'd365;value2=32'd366;
#400 value1=32'd382;value2=32'd384;
#400 value1=32'd406;value2=32'd442;
#400 value1=32'd490;value2=32'd492;
#400 value1=32'd72;value2=32'd132;
#400 value1=32'd163;value2=32'd214;
#400 value1=32'd276;value2=32'd280;
#400 value1=32'd345;value2=32'd354;
#400 value1=32'd360;value2=32'd361;
#400 value1=32'd365;value2=32'd366;
#400 value1=32'd386;value2=32'd388;
#400 value1=32'd407;value2=32'd443;
#400 value1=32'd494;value2=32'd496;
#400 value1=32'd73;value2=32'd164;
#400 value1=32'd215;value2=32'd281;
#400 value1=32'd346;value2=32'd350;
#400 value1=32'd355;value2=32'd359;
#400 value1=32'd360;value2=32'd364;
#400 value1=32'd365;value2=32'd389;
#400 value1=32'd391;value2=32'd408;
#400 value1=32'd444;value2=32'd499;
#400 value1=32'd74;value2=32'd165;
#400 value1=32'd216;value2=32'd282;
#400 value1=32'd341;value2=32'd347;
#400 value1=32'd356;value2=32'd359;
#400 value1=32'd360;value2=32'd363;
#400 value1=32'd366;value2=32'd393;
#400 value1=32'd409;value2=32'd445;
#400 value1=32'd498;value2=32'd501;
#400 value1=32'd75;value2=32'd166;
#400 value1=32'd217;value2=32'd283;
#400 value1=32'd348;value2=32'd350;
#400 value1=32'd357;value2=32'd361;
#400 value1=32'd362;value2=32'd363;
#400 value1=32'd366;value2=32'd392;
#400 value1=32'd394;value2=32'd410;
#400 value1=32'd446;value2=32'd499;
#400 value1=32'd76;value2=32'd167;
#400 value1=32'd218;value2=32'd284;
#400 value1=32'd341;value2=32'd349;
#400 value1=32'd358;value2=32'd361;
#400 value1=32'd362;value2=32'd364;
#400 value1=32'd365;value2=32'd393;
#400 value1=32'd411;value2=32'd447;
#400 value1=32'd500;value2=32'd503;
#400 value1=32'd43;value2=32'd77;
#400 value1=32'd133;value2=32'd168;
#400 value1=32'd212;value2=32'd277;
#400 value1=32'd369;value2=32'd370;
#400 value1=32'd371;value2=32'd374;
#400 value1=32'd376;value2=32'd377;
#400 value1=32'd412;value2=32'd448;
#400 value1=32'd506;value2=32'd508;
#400 value1=32'd42;value2=32'd44;
#400 value1=32'd78;value2=32'd169;
#400 value1=32'd211;value2=32'd213;
#400 value1=32'd369;value2=32'd372;
#400 value1=32'd373;value2=32'd374;
#400 value1=32'd381;value2=32'd382;
#400 value1=32'd413;value2=32'd449;
#400 value1=32'd511;value2=32'd513;
#400 value1=32'd45;value2=32'd79;
#400 value1=32'd133;value2=32'd170;
#400 value1=32'd214;value2=32'd277;
#400 value1=32'd367;value2=32'd368;
#400 value1=32'd372;value2=32'd373;
#400 value1=32'd375;value2=32'd380;
#400 value1=32'd385;value2=32'd386;
#400 value1=32'd414;value2=32'd450;
#400 value1=32'd515;value2=32'd517;
#400 value1=32'd46;value2=32'd80;
#400 value1=32'd171;value2=32'd215;
#400 value1=32'd351;value2=32'd367;
#400 value1=32'd371;value2=32'd372;
#400 value1=32'd376;value2=32'd381;
#400 value1=32'd389;value2=32'd415;
#400 value1=32'd451;value2=32'd520;
#400 value1=32'd47;value2=32'd81;
#400 value1=32'd172;value2=32'd216;
#400 value1=32'd342;value2=32'd359;
#400 value1=32'd367;value2=32'd370;
#400 value1=32'd373;value2=32'd377;
#400 value1=32'd382;value2=32'd389;
#400 value1=32'd416;value2=32'd452;
#400 value1=32'd519;value2=32'd522;
#400 value1=32'd48;value2=32'd82;
#400 value1=32'd173;value2=32'd217;
#400 value1=32'd351;value2=32'd368;
#400 value1=32'd369;value2=32'd370;
#400 value1=32'd373;value2=32'd378;
#400 value1=32'd383;value2=32'd390;
#400 value1=32'd392;value2=32'd417;
#400 value1=32'd453;value2=32'd520;
#400 value1=32'd49;value2=32'd83;
#400 value1=32'd174;value2=32'd218;
#400 value1=32'd342;value2=32'd359;
#400 value1=32'd368;value2=32'd369;
#400 value1=32'd371;value2=32'd372;
#400 value1=32'd379;value2=32'd384;
#400 value1=32'd391;value2=32'd393;
#400 value1=32'd418;value2=32'd454;
#400 value1=32'd521;value2=32'd524;
#400 value1=32'd43;value2=32'd84;
#400 value1=32'd135;value2=32'd175;
#400 value1=32'd212;value2=32'd279;
#400 value1=32'd367;value2=32'd368;
#400 value1=32'd375;value2=32'd378;
#400 value1=32'd379;value2=32'd380;
#400 value1=32'd381;value2=32'd382;
#400 value1=32'd419;value2=32'd455;
#400 value1=32'd526;value2=32'd528;
#400 value1=32'd85;value2=32'd134;
#400 value1=32'd136;value2=32'd176;
#400 value1=32'd278;value2=32'd280;
#400 value1=32'd369;value2=32'd374;
#400 value1=32'd378;value2=32'd379;
#400 value1=32'd385;value2=32'd386;
#400 value1=32'd420;value2=32'd456;
#400 value1=32'd530;value2=32'd532;
#400 value1=32'd86;value2=32'd137;
#400 value1=32'd177;value2=32'd281;
#400 value1=32'd352;value2=32'd367;
#400 value1=32'd370;value2=32'd377;
#400 value1=32'd378;value2=32'd385;
#400 value1=32'd389;value2=32'd421;
#400 value1=32'd457;value2=32'd535;
#400 value1=32'd87;value2=32'd138;
#400 value1=32'd178;value2=32'd282;
#400 value1=32'd343;value2=32'd360;
#400 value1=32'd367;value2=32'd371;
#400 value1=32'd376;value2=32'd379;
#400 value1=32'd386;value2=32'd389;
#400 value1=32'd422;value2=32'd458;
#400 value1=32'd534;value2=32'd537;
#400 value1=32'd88;value2=32'd139;
#400 value1=32'd179;value2=32'd283;
#400 value1=32'd352;value2=32'd372;
#400 value1=32'd374;value2=32'd375;
#400 value1=32'd376;value2=32'd379;
#400 value1=32'd387;value2=32'd390;
#400 value1=32'd392;value2=32'd423;
#400 value1=32'd459;value2=32'd535;
#400 value1=32'd89;value2=32'd140;
#400 value1=32'd180;value2=32'd284;
#400 value1=32'd343;value2=32'd360;
#400 value1=32'd373;value2=32'd374;
#400 value1=32'd375;value2=32'd377;
#400 value1=32'd378;value2=32'd388;
#400 value1=32'd391;value2=32'd393;
#400 value1=32'd424;value2=32'd460;
#400 value1=32'd536;value2=32'd539;
#400 value1=32'd45;value2=32'd90;
#400 value1=32'd135;value2=32'd181;
#400 value1=32'd214;value2=32'd279;
#400 value1=32'd369;value2=32'd374;
#400 value1=32'd383;value2=32'd384;
#400 value1=32'd387;value2=32'd388;
#400 value1=32'd425;value2=32'd461;
#400 value1=32'd540;value2=32'd542;
#400 value1=32'd46;value2=32'd91;
#400 value1=32'd182;value2=32'd215;
#400 value1=32'd353;value2=32'd368;
#400 value1=32'd370;value2=32'd374;
#400 value1=32'd382;value2=32'd383;
#400 value1=32'd385;value2=32'd390;
#400 value1=32'd391;value2=32'd426;
#400 value1=32'd462;value2=32'd545;
#400 value1=32'd47;value2=32'd92;
#400 value1=32'd183;value2=32'd216;
#400 value1=32'd344;value2=32'd361;
#400 value1=32'd368;value2=32'd371;
#400 value1=32'd374;value2=32'd381;
#400 value1=32'd384;value2=32'd386;
#400 value1=32'd392;value2=32'd393;
#400 value1=32'd427;value2=32'd463;
#400 value1=32'd544;value2=32'd547;
#400 value1=32'd48;value2=32'd93;
#400 value1=32'd184;value2=32'd217;
#400 value1=32'd353;value2=32'd372;
#400 value1=32'd380;value2=32'd381;
#400 value1=32'd384;value2=32'd387;
#400 value1=32'd394;value2=32'd428;
#400 value1=32'd464;value2=32'd545;
#400 value1=32'd49;value2=32'd94;
#400 value1=32'd185;value2=32'd218;
#400 value1=32'd344;value2=32'd361;
#400 value1=32'd373;value2=32'd380;
#400 value1=32'd382;value2=32'd383;
#400 value1=32'd388;value2=32'd394;
#400 value1=32'd429;value2=32'd465;
#400 value1=32'd546;value2=32'd549;
#400 value1=32'd95;value2=32'd137;
#400 value1=32'd186;value2=32'd281;
#400 value1=32'd354;value2=32'd369;
#400 value1=32'd375;value2=32'd376;
#400 value1=32'd381;value2=32'd386;
#400 value1=32'd387;value2=32'd390;
#400 value1=32'd391;value2=32'd430;
#400 value1=32'd466;value2=32'd551;
#400 value1=32'd96;value2=32'd138;
#400 value1=32'd187;value2=32'd282;
#400 value1=32'd345;value2=32'd362;
#400 value1=32'd369;value2=32'd375;
#400 value1=32'd377;value2=32'd382;
#400 value1=32'd385;value2=32'd388;
#400 value1=32'd392;value2=32'd393;
#400 value1=32'd431;value2=32'd467;
#400 value1=32'd550;value2=32'd553;
#400 value1=32'd97;value2=32'd139;
#400 value1=32'd188;value2=32'd283;
#400 value1=32'd354;value2=32'd378;
#400 value1=32'd380;value2=32'd383;
#400 value1=32'd385;value2=32'd388;
#400 value1=32'd394;value2=32'd432;
#400 value1=32'd468;value2=32'd551;
#400 value1=32'd98;value2=32'd140;
#400 value1=32'd189;value2=32'd284;
#400 value1=32'd345;value2=32'd362;
#400 value1=32'd379;value2=32'd380;
#400 value1=32'd384;value2=32'd386;
#400 value1=32'd387;value2=32'd394;
#400 value1=32'd433;value2=32'd469;
#400 value1=32'd552;value2=32'd555;
#400 value1=32'd99;value2=32'd190;
#400 value1=32'd346;value2=32'd356;
#400 value1=32'd363;value2=32'd370;
#400 value1=32'd371;value2=32'd376;
#400 value1=32'd377;value2=32'd391;
#400 value1=32'd392;value2=32'd434;
#400 value1=32'd470;value2=32'd556;
#400 value1=32'd100;value2=32'd191;
#400 value1=32'd355;value2=32'd357;
#400 value1=32'd372;value2=32'd378;
#400 value1=32'd381;value2=32'd385;
#400 value1=32'd391;value2=32'd392;
#400 value1=32'd435;value2=32'd471;
#400 value1=32'd101;value2=32'd192;
#400 value1=32'd346;value2=32'd358;
#400 value1=32'd363;value2=32'd373;
#400 value1=32'd379;value2=32'd381;
#400 value1=32'd385;value2=32'd389;
#400 value1=32'd390;value2=32'd393;
#400 value1=32'd394;value2=32'd436;
#400 value1=32'd472;value2=32'd558;
#400 value1=32'd102;value2=32'd193;
#400 value1=32'd348;value2=32'd356;
#400 value1=32'd365;value2=32'd372;
#400 value1=32'd378;value2=32'd382;
#400 value1=32'd386;value2=32'd389;
#400 value1=32'd390;value2=32'd393;
#400 value1=32'd394;value2=32'd437;
#400 value1=32'd473;value2=32'd556;
#400 value1=32'd103;value2=32'd194;
#400 value1=32'd347;value2=32'd349;
#400 value1=32'd364;value2=32'd366;
#400 value1=32'd373;value2=32'd379;
#400 value1=32'd382;value2=32'd386;
#400 value1=32'd391;value2=32'd392;
#400 value1=32'd438;value2=32'd474;
#400 value1=32'd557;value2=32'd559;
#400 value1=32'd104;value2=32'd195;
#400 value1=32'd348;value2=32'd358;
#400 value1=32'd365;value2=32'd383;
#400 value1=32'd384;value2=32'd387;
#400 value1=32'd388;value2=32'd391;
#400 value1=32'd392;value2=32'd439;
#400 value1=32'd475;value2=32'd558;
#400 value1=32'd60;value2=32'd151;
#400 value1=32'd219;value2=32'd220;
#400 value1=32'd285;value2=32'd286;
#400 value1=32'd341;value2=32'd350;
#400 value1=32'd401;value2=32'd403;
#400 value1=32'd408;value2=32'd410;
#400 value1=32'd445;value2=32'd447;
#400 value1=32'd50;value2=32'd61;
#400 value1=32'd152;value2=32'd219;
#400 value1=32'd221;value2=32'd287;
#400 value1=32'd342;value2=32'd351;
#400 value1=32'd397;value2=32'd398;
#400 value1=32'd400;value2=32'd401;
#400 value1=32'd404;value2=32'd415;
#400 value1=32'd417;value2=32'd440;
#400 value1=32'd452;value2=32'd454;
#400 value1=32'd62;value2=32'd141;
#400 value1=32'd153;value2=32'd222;
#400 value1=32'd285;value2=32'd288;
#400 value1=32'd343;value2=32'd352;
#400 value1=32'd396;value2=32'd399;
#400 value1=32'd400;value2=32'd401;
#400 value1=32'd405;value2=32'd421;
#400 value1=32'd423;value2=32'd441;
#400 value1=32'd458;value2=32'd460;
#400 value1=32'd50;value2=32'd63;
#400 value1=32'd154;value2=32'd219;
#400 value1=32'd223;value2=32'd289;
#400 value1=32'd344;value2=32'd353;
#400 value1=32'd396;value2=32'd399;
#400 value1=32'd402;value2=32'd403;
#400 value1=32'd406;value2=32'd426;
#400 value1=32'd428;value2=32'd442;
#400 value1=32'd463;value2=32'd465;
#400 value1=32'd64;value2=32'd141;
#400 value1=32'd155;value2=32'd224;
#400 value1=32'd285;value2=32'd290;
#400 value1=32'd345;value2=32'd354;
#400 value1=32'd397;value2=32'd398;
#400 value1=32'd402;value2=32'd403;
#400 value1=32'd407;value2=32'd430;
#400 value1=32'd432;value2=32'd443;
#400 value1=32'd467;value2=32'd469;
#400 value1=32'd65;value2=32'd156;
#400 value1=32'd225;value2=32'd291;
#400 value1=32'd340;value2=32'd346;
#400 value1=32'd355;value2=32'd396;
#400 value1=32'd397;value2=32'd401;
#400 value1=32'd402;value2=32'd408;
#400 value1=32'd435;value2=32'd444;
#400 value1=32'd470;value2=32'd472;
#400 value1=32'd66;value2=32'd157;
#400 value1=32'd226;value2=32'd292;
#400 value1=32'd347;value2=32'd356;
#400 value1=32'd395;value2=32'd396;
#400 value1=32'd397;value2=32'd400;
#400 value1=32'd403;value2=32'd409;
#400 value1=32'd434;value2=32'd437;
#400 value1=32'd445;value2=32'd474;
#400 value1=32'd67;value2=32'd158;
#400 value1=32'd227;value2=32'd293;
#400 value1=32'd340;value2=32'd348;
#400 value1=32'd357;value2=32'd398;
#400 value1=32'd399;value2=32'd400;
#400 value1=32'd403;value2=32'd410;
#400 value1=32'd435;value2=32'd446;
#400 value1=32'd473;value2=32'd475;
#400 value1=32'd68;value2=32'd159;
#400 value1=32'd228;value2=32'd294;
#400 value1=32'd349;value2=32'd358;
#400 value1=32'd395;value2=32'd398;
#400 value1=32'd399;value2=32'd401;
#400 value1=32'd402;value2=32'd411;
#400 value1=32'd436;value2=32'd439;
#400 value1=32'd447;value2=32'd474;
#400 value1=32'd51;value2=32'd69;
#400 value1=32'd160;value2=32'd220;
#400 value1=32'd221;value2=32'd287;
#400 value1=32'd359;value2=32'd396;
#400 value1=32'd405;value2=32'd406;
#400 value1=32'd408;value2=32'd409;
#400 value1=32'd416;value2=32'd418;
#400 value1=32'd480;value2=32'd482;
#400 value1=32'd70;value2=32'd142;
#400 value1=32'd161;value2=32'd222;
#400 value1=32'd286;value2=32'd288;
#400 value1=32'd360;value2=32'd397;
#400 value1=32'd404;value2=32'd407;
#400 value1=32'd408;value2=32'd409;
#400 value1=32'd422;value2=32'd424;
#400 value1=32'd486;value2=32'd488;
#400 value1=32'd51;value2=32'd71;
#400 value1=32'd162;value2=32'd220;
#400 value1=32'd223;value2=32'd289;
#400 value1=32'd361;value2=32'd398;
#400 value1=32'd404;value2=32'd407;
#400 value1=32'd410;value2=32'd411;
#400 value1=32'd427;value2=32'd429;
#400 value1=32'd491;value2=32'd493;
#400 value1=32'd72;value2=32'd142;
#400 value1=32'd163;value2=32'd224;
#400 value1=32'd286;value2=32'd290;
#400 value1=32'd362;value2=32'd399;
#400 value1=32'd405;value2=32'd406;
#400 value1=32'd410;value2=32'd411;
#400 value1=32'd431;value2=32'd433;
#400 value1=32'd495;value2=32'd497;
#400 value1=32'd73;value2=32'd164;
#400 value1=32'd225;value2=32'd291;
#400 value1=32'd341;value2=32'd363;
#400 value1=32'd395;value2=32'd400;
#400 value1=32'd404;value2=32'd405;
#400 value1=32'd409;value2=32'd410;
#400 value1=32'd434;value2=32'd436;
#400 value1=32'd498;value2=32'd500;
#400 value1=32'd74;value2=32'd165;
#400 value1=32'd226;value2=32'd292;
#400 value1=32'd364;value2=32'd401;
#400 value1=32'd404;value2=32'd405;
#400 value1=32'd408;value2=32'd411;
#400 value1=32'd438;value2=32'd502;
#400 value1=32'd75;value2=32'd166;
#400 value1=32'd227;value2=32'd293;
#400 value1=32'd341;value2=32'd365;
#400 value1=32'd395;value2=32'd402;
#400 value1=32'd406;value2=32'd407;
#400 value1=32'd408;value2=32'd411;
#400 value1=32'd437;value2=32'd439;
#400 value1=32'd501;value2=32'd503;
#400 value1=32'd76;value2=32'd167;
#400 value1=32'd228;value2=32'd294;
#400 value1=32'd366;value2=32'd403;
#400 value1=32'd406;value2=32'd407;
#400 value1=32'd409;value2=32'd410;
#400 value1=32'd438;value2=32'd502;
#400 value1=32'd53;value2=32'd77;
#400 value1=32'd143;value2=32'd168;
#400 value1=32'd222;value2=32'd287;
#400 value1=32'd367;value2=32'd414;
#400 value1=32'd415;value2=32'd416;
#400 value1=32'd419;value2=32'd421;
#400 value1=32'd422;value2=32'd476;
#400 value1=32'd507;value2=32'd509;
#400 value1=32'd52;value2=32'd54;
#400 value1=32'd78;value2=32'd169;
#400 value1=32'd221;value2=32'd223;
#400 value1=32'd368;value2=32'd414;
#400 value1=32'd417;value2=32'd418;
#400 value1=32'd419;value2=32'd426;
#400 value1=32'd427;value2=32'd477;
#400 value1=32'd512;value2=32'd514;
#400 value1=32'd55;value2=32'd79;
#400 value1=32'd143;value2=32'd170;
#400 value1=32'd224;value2=32'd287;
#400 value1=32'd369;value2=32'd412;
#400 value1=32'd413;value2=32'd417;
#400 value1=32'd418;value2=32'd420;
#400 value1=32'd425;value2=32'd430;
#400 value1=32'd431;value2=32'd478;
#400 value1=32'd516;value2=32'd518;
#400 value1=32'd56;value2=32'd80;
#400 value1=32'd171;value2=32'd225;
#400 value1=32'd342;value2=32'd370;
#400 value1=32'd396;value2=32'd412;
#400 value1=32'd416;value2=32'd417;
#400 value1=32'd421;value2=32'd426;
#400 value1=32'd434;value2=32'd479;
#400 value1=32'd519;value2=32'd521;
#400 value1=32'd57;value2=32'd81;
#400 value1=32'd172;value2=32'd226;
#400 value1=32'd371;value2=32'd404;
#400 value1=32'd412;value2=32'd415;
#400 value1=32'd418;value2=32'd422;
#400 value1=32'd427;value2=32'd434;
#400 value1=32'd480;value2=32'd523;
#400 value1=32'd58;value2=32'd82;
#400 value1=32'd173;value2=32'd227;
#400 value1=32'd342;value2=32'd372;
#400 value1=32'd396;value2=32'd413;
#400 value1=32'd414;value2=32'd415;
#400 value1=32'd418;value2=32'd423;
#400 value1=32'd428;value2=32'd435;
#400 value1=32'd437;value2=32'd481;
#400 value1=32'd522;value2=32'd524;
#400 value1=32'd59;value2=32'd83;
#400 value1=32'd174;value2=32'd228;
#400 value1=32'd373;value2=32'd404;
#400 value1=32'd413;value2=32'd414;
#400 value1=32'd416;value2=32'd417;
#400 value1=32'd424;value2=32'd429;
#400 value1=32'd436;value2=32'd438;
#400 value1=32'd482;value2=32'd523;
#400 value1=32'd53;value2=32'd84;
#400 value1=32'd145;value2=32'd175;
#400 value1=32'd222;value2=32'd289;
#400 value1=32'd374;value2=32'd412;
#400 value1=32'd413;value2=32'd420;
#400 value1=32'd423;value2=32'd424;
#400 value1=32'd425;value2=32'd426;
#400 value1=32'd427;value2=32'd483;
#400 value1=32'd527;value2=32'd529;
#400 value1=32'd85;value2=32'd144;
#400 value1=32'd146;value2=32'd176;
#400 value1=32'd288;value2=32'd290;
#400 value1=32'd375;value2=32'd414;
#400 value1=32'd419;value2=32'd423;
#400 value1=32'd424;value2=32'd430;
#400 value1=32'd431;value2=32'd484;
#400 value1=32'd531;value2=32'd533;
#400 value1=32'd86;value2=32'd147;
#400 value1=32'd177;value2=32'd291;
#400 value1=32'd343;value2=32'd376;
#400 value1=32'd397;value2=32'd412;
#400 value1=32'd415;value2=32'd422;
#400 value1=32'd423;value2=32'd430;
#400 value1=32'd434;value2=32'd485;
#400 value1=32'd534;value2=32'd536;
#400 value1=32'd87;value2=32'd148;
#400 value1=32'd178;value2=32'd292;
#400 value1=32'd377;value2=32'd405;
#400 value1=32'd412;value2=32'd416;
#400 value1=32'd421;value2=32'd424;
#400 value1=32'd431;value2=32'd434;
#400 value1=32'd486;value2=32'd538;
#400 value1=32'd88;value2=32'd149;
#400 value1=32'd179;value2=32'd293;
#400 value1=32'd343;value2=32'd378;
#400 value1=32'd397;value2=32'd417;
#400 value1=32'd419;value2=32'd420;
#400 value1=32'd421;value2=32'd424;
#400 value1=32'd432;value2=32'd435;
#400 value1=32'd437;value2=32'd487;
#400 value1=32'd537;value2=32'd539;
#400 value1=32'd89;value2=32'd150;
#400 value1=32'd180;value2=32'd294;
#400 value1=32'd379;value2=32'd405;
#400 value1=32'd418;value2=32'd419;
#400 value1=32'd420;value2=32'd422;
#400 value1=32'd423;value2=32'd433;
#400 value1=32'd436;value2=32'd438;
#400 value1=32'd488;value2=32'd538;
#400 value1=32'd55;value2=32'd90;
#400 value1=32'd145;value2=32'd181;
#400 value1=32'd224;value2=32'd289;
#400 value1=32'd380;value2=32'd414;
#400 value1=32'd419;value2=32'd428;
#400 value1=32'd429;value2=32'd432;
#400 value1=32'd433;value2=32'd489;
#400 value1=32'd541;value2=32'd543;
#400 value1=32'd56;value2=32'd91;
#400 value1=32'd182;value2=32'd225;
#400 value1=32'd344;value2=32'd381;
#400 value1=32'd398;value2=32'd413;
#400 value1=32'd415;value2=32'd419;
#400 value1=32'd427;value2=32'd428;
#400 value1=32'd430;value2=32'd435;
#400 value1=32'd436;value2=32'd490;
#400 value1=32'd544;value2=32'd546;
#400 value1=32'd57;value2=32'd92;
#400 value1=32'd183;value2=32'd226;
#400 value1=32'd382;value2=32'd406;
#400 value1=32'd413;value2=32'd416;
#400 value1=32'd419;value2=32'd426;
#400 value1=32'd429;value2=32'd431;
#400 value1=32'd437;value2=32'd438;
#400 value1=32'd491;value2=32'd548;
#400 value1=32'd58;value2=32'd93;
#400 value1=32'd184;value2=32'd227;
#400 value1=32'd344;value2=32'd383;
#400 value1=32'd398;value2=32'd417;
#400 value1=32'd425;value2=32'd426;
#400 value1=32'd429;value2=32'd432;
#400 value1=32'd439;value2=32'd492;
#400 value1=32'd547;value2=32'd549;
#400 value1=32'd59;value2=32'd94;
#400 value1=32'd185;value2=32'd228;
#400 value1=32'd384;value2=32'd406;
#400 value1=32'd418;value2=32'd425;
#400 value1=32'd427;value2=32'd428;
#400 value1=32'd433;value2=32'd439;
#400 value1=32'd493;value2=32'd548;
#400 value1=32'd95;value2=32'd147;
#400 value1=32'd186;value2=32'd291;
#400 value1=32'd345;value2=32'd385;
#400 value1=32'd399;value2=32'd414;
#400 value1=32'd420;value2=32'd421;
#400 value1=32'd426;value2=32'd431;
#400 value1=32'd432;value2=32'd435;
#400 value1=32'd436;value2=32'd494;
#400 value1=32'd550;value2=32'd552;
#400 value1=32'd96;value2=32'd148;
#400 value1=32'd187;value2=32'd292;
#400 value1=32'd386;value2=32'd407;
#400 value1=32'd414;value2=32'd420;
#400 value1=32'd422;value2=32'd427;
#400 value1=32'd430;value2=32'd433;
#400 value1=32'd437;value2=32'd438;
#400 value1=32'd495;value2=32'd554;
#400 value1=32'd97;value2=32'd149;
#400 value1=32'd188;value2=32'd293;
#400 value1=32'd345;value2=32'd387;
#400 value1=32'd399;value2=32'd423;
#400 value1=32'd425;value2=32'd428;
#400 value1=32'd430;value2=32'd433;
#400 value1=32'd439;value2=32'd496;
#400 value1=32'd553;value2=32'd555;
#400 value1=32'd98;value2=32'd150;
#400 value1=32'd189;value2=32'd294;
#400 value1=32'd388;value2=32'd407;
#400 value1=32'd424;value2=32'd425;
#400 value1=32'd429;value2=32'd431;
#400 value1=32'd432;value2=32'd439;
#400 value1=32'd497;value2=32'd554;
#400 value1=32'd99;value2=32'd190;
#400 value1=32'd347;value2=32'd389;
#400 value1=32'd401;value2=32'd408;
#400 value1=32'd415;value2=32'd416;
#400 value1=32'd421;value2=32'd422;
#400 value1=32'd436;value2=32'd437;
#400 value1=32'd498;value2=32'd557;
#400 value1=32'd100;value2=32'd191;
#400 value1=32'd346;value2=32'd348;
#400 value1=32'd390;value2=32'd400;
#400 value1=32'd402;value2=32'd417;
#400 value1=32'd423;value2=32'd426;
#400 value1=32'd430;value2=32'd436;
#400 value1=32'd437;value2=32'd499;
#400 value1=32'd556;value2=32'd558;
#400 value1=32'd101;value2=32'd192;
#400 value1=32'd349;value2=32'd391;
#400 value1=32'd403;value2=32'd408;
#400 value1=32'd418;value2=32'd424;
#400 value1=32'd426;value2=32'd430;
#400 value1=32'd434;value2=32'd435;
#400 value1=32'd438;value2=32'd439;
#400 value1=32'd500;value2=32'd557;
#400 value1=32'd102;value2=32'd193;
#400 value1=32'd347;value2=32'd392;
#400 value1=32'd401;value2=32'd410;
#400 value1=32'd417;value2=32'd423;
#400 value1=32'd427;value2=32'd431;
#400 value1=32'd434;value2=32'd435;
#400 value1=32'd438;value2=32'd439;
#400 value1=32'd501;value2=32'd559;
#400 value1=32'd103;value2=32'd194;
#400 value1=32'd393;value2=32'd409;
#400 value1=32'd411;value2=32'd418;
#400 value1=32'd424;value2=32'd427;
#400 value1=32'd431;value2=32'd436;
#400 value1=32'd437;value2=32'd502;
#400 value1=32'd104;value2=32'd195;
#400 value1=32'd349;value2=32'd394;
#400 value1=32'd403;value2=32'd410;
#400 value1=32'd428;value2=32'd429;
#400 value1=32'd432;value2=32'd433;
#400 value1=32'd436;value2=32'd437;
#400 value1=32'd503;value2=32'd559;
#400 value1=32'd60;value2=32'd229;
#400 value1=32'd230;value2=32'd238;
#400 value1=32'd296;value2=32'd304;
#400 value1=32'd359;value2=32'd396;
#400 value1=32'd441;value2=32'd442;
#400 value1=32'd444;value2=32'd445;
#400 value1=32'd452;value2=32'd454;
#400 value1=32'd479;value2=32'd481;
#400 value1=32'd151;value2=32'd231;
#400 value1=32'd239;value2=32'd295;
#400 value1=32'd297;value2=32'd305;
#400 value1=32'd360;value2=32'd397;
#400 value1=32'd440;value2=32'd443;
#400 value1=32'd444;value2=32'd445;
#400 value1=32'd458;value2=32'd460;
#400 value1=32'd485;value2=32'd487;
#400 value1=32'd60;value2=32'd229;
#400 value1=32'd232;value2=32'd240;
#400 value1=32'd298;value2=32'd306;
#400 value1=32'd361;value2=32'd398;
#400 value1=32'd440;value2=32'd443;
#400 value1=32'd446;value2=32'd447;
#400 value1=32'd463;value2=32'd465;
#400 value1=32'd490;value2=32'd492;
#400 value1=32'd151;value2=32'd233;
#400 value1=32'd241;value2=32'd295;
#400 value1=32'd299;value2=32'd307;
#400 value1=32'd362;value2=32'd399;
#400 value1=32'd441;value2=32'd442;
#400 value1=32'd446;value2=32'd447;
#400 value1=32'd467;value2=32'd469;
#400 value1=32'd494;value2=32'd496;
#400 value1=32'd234;value2=32'd242;
#400 value1=32'd300;value2=32'd308;
#400 value1=32'd350;value2=32'd363;
#400 value1=32'd400;value2=32'd440;
#400 value1=32'd441;value2=32'd445;
#400 value1=32'd446;value2=32'd470;
#400 value1=32'd472;value2=32'd499;
#400 value1=32'd235;value2=32'd243;
#400 value1=32'd301;value2=32'd309;
#400 value1=32'd364;value2=32'd395;
#400 value1=32'd401;value2=32'd440;
#400 value1=32'd441;value2=32'd444;
#400 value1=32'd447;value2=32'd474;
#400 value1=32'd498;value2=32'd501;
#400 value1=32'd236;value2=32'd244;
#400 value1=32'd302;value2=32'd310;
#400 value1=32'd350;value2=32'd365;
#400 value1=32'd402;value2=32'd442;
#400 value1=32'd443;value2=32'd444;
#400 value1=32'd447;value2=32'd473;
#400 value1=32'd475;value2=32'd499;
#400 value1=32'd237;value2=32'd245;
#400 value1=32'd303;value2=32'd311;
#400 value1=32'd366;value2=32'd395;
#400 value1=32'd403;value2=32'd442;
#400 value1=32'd443;value2=32'd445;
#400 value1=32'd446;value2=32'd474;
#400 value1=32'd500;value2=32'd503;
#400 value1=32'd62;value2=32'd152;
#400 value1=32'd231;value2=32'd246;
#400 value1=32'd296;value2=32'd312;
#400 value1=32'd367;value2=32'd450;
#400 value1=32'd451;value2=32'd452;
#400 value1=32'd455;value2=32'd457;
#400 value1=32'd458;value2=32'd476;
#400 value1=32'd506;value2=32'd508;
#400 value1=32'd61;value2=32'd63;
#400 value1=32'd230;value2=32'd232;
#400 value1=32'd247;value2=32'd313;
#400 value1=32'd368;value2=32'd450;
#400 value1=32'd453;value2=32'd454;
#400 value1=32'd455;value2=32'd462;
#400 value1=32'd463;value2=32'd477;
#400 value1=32'd511;value2=32'd513;
#400 value1=32'd64;value2=32'd152;
#400 value1=32'd233;value2=32'd248;
#400 value1=32'd296;value2=32'd314;
#400 value1=32'd369;value2=32'd448;
#400 value1=32'd449;value2=32'd453;
#400 value1=32'd454;value2=32'd456;
#400 value1=32'd461;value2=32'd466;
#400 value1=32'd467;value2=32'd478;
#400 value1=32'd515;value2=32'd517;
#400 value1=32'd65;value2=32'd234;
#400 value1=32'd249;value2=32'd315;
#400 value1=32'd351;value2=32'd370;
#400 value1=32'd448;value2=32'd452;
#400 value1=32'd453;value2=32'd457;
#400 value1=32'd462;value2=32'd470;
#400 value1=32'd479;value2=32'd520;
#400 value1=32'd66;value2=32'd235;
#400 value1=32'd250;value2=32'd316;
#400 value1=32'd371;value2=32'd396;
#400 value1=32'd440;value2=32'd448;
#400 value1=32'd451;value2=32'd454;
#400 value1=32'd458;value2=32'd463;
#400 value1=32'd470;value2=32'd480;
#400 value1=32'd519;value2=32'd522;
#400 value1=32'd67;value2=32'd236;
#400 value1=32'd251;value2=32'd317;
#400 value1=32'd351;value2=32'd372;
#400 value1=32'd449;value2=32'd450;
#400 value1=32'd451;value2=32'd454;
#400 value1=32'd459;value2=32'd464;
#400 value1=32'd471;value2=32'd473;
#400 value1=32'd481;value2=32'd520;
#400 value1=32'd68;value2=32'd237;
#400 value1=32'd252;value2=32'd318;
#400 value1=32'd373;value2=32'd396;
#400 value1=32'd440;value2=32'd449;
#400 value1=32'd450;value2=32'd452;
#400 value1=32'd453;value2=32'd460;
#400 value1=32'd465;value2=32'd472;
#400 value1=32'd474;value2=32'd482;
#400 value1=32'd521;value2=32'd524;
#400 value1=32'd62;value2=32'd154;
#400 value1=32'd231;value2=32'd253;
#400 value1=32'd298;value2=32'd319;
#400 value1=32'd374;value2=32'd448;
#400 value1=32'd449;value2=32'd456;
#400 value1=32'd459;value2=32'd460;
#400 value1=32'd461;value2=32'd462;
#400 value1=32'd463;value2=32'd483;
#400 value1=32'd526;value2=32'd528;
#400 value1=32'd153;value2=32'd155;
#400 value1=32'd254;value2=32'd297;
#400 value1=32'd299;value2=32'd320;
#400 value1=32'd375;value2=32'd450;
#400 value1=32'd455;value2=32'd459;
#400 value1=32'd460;value2=32'd466;
#400 value1=32'd467;value2=32'd484;
#400 value1=32'd530;value2=32'd532;
#400 value1=32'd156;value2=32'd255;
#400 value1=32'd300;value2=32'd321;
#400 value1=32'd352;value2=32'd376;
#400 value1=32'd448;value2=32'd451;
#400 value1=32'd458;value2=32'd459;
#400 value1=32'd466;value2=32'd470;
#400 value1=32'd485;value2=32'd535;
#400 value1=32'd157;value2=32'd256;
#400 value1=32'd301;value2=32'd322;
#400 value1=32'd377;value2=32'd397;
#400 value1=32'd441;value2=32'd448;
#400 value1=32'd452;value2=32'd457;
#400 value1=32'd460;value2=32'd467;
#400 value1=32'd470;value2=32'd486;
#400 value1=32'd534;value2=32'd537;
#400 value1=32'd158;value2=32'd257;
#400 value1=32'd302;value2=32'd323;
#400 value1=32'd352;value2=32'd378;
#400 value1=32'd453;value2=32'd455;
#400 value1=32'd456;value2=32'd457;
#400 value1=32'd460;value2=32'd468;
#400 value1=32'd471;value2=32'd473;
#400 value1=32'd487;value2=32'd535;
#400 value1=32'd159;value2=32'd258;
#400 value1=32'd303;value2=32'd324;
#400 value1=32'd379;value2=32'd397;
#400 value1=32'd441;value2=32'd454;
#400 value1=32'd455;value2=32'd456;
#400 value1=32'd458;value2=32'd459;
#400 value1=32'd469;value2=32'd472;
#400 value1=32'd474;value2=32'd488;
#400 value1=32'd536;value2=32'd539;
#400 value1=32'd64;value2=32'd154;
#400 value1=32'd233;value2=32'd259;
#400 value1=32'd298;value2=32'd325;
#400 value1=32'd380;value2=32'd450;
#400 value1=32'd455;value2=32'd464;
#400 value1=32'd465;value2=32'd468;
#400 value1=32'd469;value2=32'd489;
#400 value1=32'd540;value2=32'd542;
#400 value1=32'd65;value2=32'd234;
#400 value1=32'd260;value2=32'd326;
#400 value1=32'd353;value2=32'd381;
#400 value1=32'd449;value2=32'd451;
#400 value1=32'd455;value2=32'd463;
#400 value1=32'd464;value2=32'd466;
#400 value1=32'd471;value2=32'd472;
#400 value1=32'd490;value2=32'd545;
#400 value1=32'd66;value2=32'd235;
#400 value1=32'd261;value2=32'd327;
#400 value1=32'd382;value2=32'd398;
#400 value1=32'd442;value2=32'd449;
#400 value1=32'd452;value2=32'd455;
#400 value1=32'd462;value2=32'd465;
#400 value1=32'd467;value2=32'd473;
#400 value1=32'd474;value2=32'd491;
#400 value1=32'd544;value2=32'd547;
#400 value1=32'd67;value2=32'd236;
#400 value1=32'd262;value2=32'd328;
#400 value1=32'd353;value2=32'd383;
#400 value1=32'd453;value2=32'd461;
#400 value1=32'd462;value2=32'd465;
#400 value1=32'd468;value2=32'd475;
#400 value1=32'd492;value2=32'd545;
#400 value1=32'd68;value2=32'd237;
#400 value1=32'd263;value2=32'd329;
#400 value1=32'd384;value2=32'd398;
#400 value1=32'd442;value2=32'd454;
#400 value1=32'd461;value2=32'd463;
#400 value1=32'd464;value2=32'd469;
#400 value1=32'd475;value2=32'd493;
#400 value1=32'd546;value2=32'd549;
#400 value1=32'd156;value2=32'd264;
#400 value1=32'd300;value2=32'd330;
#400 value1=32'd354;value2=32'd385;
#400 value1=32'd450;value2=32'd456;
#400 value1=32'd457;value2=32'd462;
#400 value1=32'd467;value2=32'd468;
#400 value1=32'd471;value2=32'd472;
#400 value1=32'd494;value2=32'd551;
#400 value1=32'd157;value2=32'd265;
#400 value1=32'd301;value2=32'd331;
#400 value1=32'd386;value2=32'd399;
#400 value1=32'd443;value2=32'd450;
#400 value1=32'd456;value2=32'd458;
#400 value1=32'd463;value2=32'd466;
#400 value1=32'd469;value2=32'd473;
#400 value1=32'd474;value2=32'd495;
#400 value1=32'd550;value2=32'd553;
#400 value1=32'd158;value2=32'd266;
#400 value1=32'd302;value2=32'd332;
#400 value1=32'd354;value2=32'd387;
#400 value1=32'd459;value2=32'd461;
#400 value1=32'd464;value2=32'd466;
#400 value1=32'd469;value2=32'd475;
#400 value1=32'd496;value2=32'd551;
#400 value1=32'd159;value2=32'd267;
#400 value1=32'd303;value2=32'd333;
#400 value1=32'd388;value2=32'd399;
#400 value1=32'd443;value2=32'd460;
#400 value1=32'd461;value2=32'd465;
#400 value1=32'd467;value2=32'd468;
#400 value1=32'd475;value2=32'd497;
#400 value1=32'd552;value2=32'd555;
#400 value1=32'd268;value2=32'd334;
#400 value1=32'd356;value2=32'd389;
#400 value1=32'd400;value2=32'd444;
#400 value1=32'd451;value2=32'd452;
#400 value1=32'd457;value2=32'd458;
#400 value1=32'd472;value2=32'd473;
#400 value1=32'd498;value2=32'd556;
#400 value1=32'd269;value2=32'd335;
#400 value1=32'd355;value2=32'd357;
#400 value1=32'd390;value2=32'd453;
#400 value1=32'd459;value2=32'd462;
#400 value1=32'd466;value2=32'd472;
#400 value1=32'd473;value2=32'd499;
#400 value1=32'd270;value2=32'd336;
#400 value1=32'd358;value2=32'd391;
#400 value1=32'd400;value2=32'd444;
#400 value1=32'd454;value2=32'd460;
#400 value1=32'd462;value2=32'd466;
#400 value1=32'd470;value2=32'd471;
#400 value1=32'd474;value2=32'd475;
#400 value1=32'd500;value2=32'd558;
#400 value1=32'd271;value2=32'd337;
#400 value1=32'd356;value2=32'd392;
#400 value1=32'd402;value2=32'd446;
#400 value1=32'd453;value2=32'd459;
#400 value1=32'd463;value2=32'd467;
#400 value1=32'd470;value2=32'd471;
#400 value1=32'd474;value2=32'd475;
#400 value1=32'd501;value2=32'd556;
#400 value1=32'd272;value2=32'd338;
#400 value1=32'd393;value2=32'd401;
#400 value1=32'd403;value2=32'd445;
#400 value1=32'd447;value2=32'd454;
#400 value1=32'd460;value2=32'd463;
#400 value1=32'd467;value2=32'd472;
#400 value1=32'd473;value2=32'd502;
#400 value1=32'd557;value2=32'd559;
#400 value1=32'd273;value2=32'd339;
#400 value1=32'd358;value2=32'd394;
#400 value1=32'd402;value2=32'd446;
#400 value1=32'd464;value2=32'd465;
#400 value1=32'd468;value2=32'd469;
#400 value1=32'd472;value2=32'd473;
#400 value1=32'd503;value2=32'd558;
#400 value1=32'd70;value2=32'd160;
#400 value1=32'd239;value2=32'd246;
#400 value1=32'd304;value2=32'd312;
#400 value1=32'd412;value2=32'd448;
#400 value1=32'd478;value2=32'd479;
#400 value1=32'd480;value2=32'd483;
#400 value1=32'd485;value2=32'd486;
#400 value1=32'd507;value2=32'd509;
#400 value1=32'd69;value2=32'd71;
#400 value1=32'd238;value2=32'd240;
#400 value1=32'd247;value2=32'd313;
#400 value1=32'd413;value2=32'd449;
#400 value1=32'd478;value2=32'd481;
#400 value1=32'd482;value2=32'd483;
#400 value1=32'd490;value2=32'd491;
#400 value1=32'd512;value2=32'd514;
#400 value1=32'd72;value2=32'd160;
#400 value1=32'd241;value2=32'd248;
#400 value1=32'd304;value2=32'd314;
#400 value1=32'd414;value2=32'd450;
#400 value1=32'd476;value2=32'd477;
#400 value1=32'd481;value2=32'd482;
#400 value1=32'd484;value2=32'd489;
#400 value1=32'd494;value2=32'd495;
#400 value1=32'd516;value2=32'd518;
#400 value1=32'd73;value2=32'd242;
#400 value1=32'd249;value2=32'd315;
#400 value1=32'd359;value2=32'd415;
#400 value1=32'd440;value2=32'd451;
#400 value1=32'd476;value2=32'd480;
#400 value1=32'd481;value2=32'd485;
#400 value1=32'd490;value2=32'd498;
#400 value1=32'd519;value2=32'd521;
#400 value1=32'd74;value2=32'd243;
#400 value1=32'd250;value2=32'd316;
#400 value1=32'd404;value2=32'd416;
#400 value1=32'd452;value2=32'd476;
#400 value1=32'd479;value2=32'd482;
#400 value1=32'd486;value2=32'd491;
#400 value1=32'd498;value2=32'd523;
#400 value1=32'd75;value2=32'd244;
#400 value1=32'd251;value2=32'd317;
#400 value1=32'd359;value2=32'd417;
#400 value1=32'd440;value2=32'd453;
#400 value1=32'd477;value2=32'd478;
#400 value1=32'd479;value2=32'd482;
#400 value1=32'd487;value2=32'd492;
#400 value1=32'd499;value2=32'd501;
#400 value1=32'd522;value2=32'd524;
#400 value1=32'd76;value2=32'd245;
#400 value1=32'd252;value2=32'd318;
#400 value1=32'd404;value2=32'd418;
#400 value1=32'd454;value2=32'd477;
#400 value1=32'd478;value2=32'd480;
#400 value1=32'd481;value2=32'd488;
#400 value1=32'd493;value2=32'd500;
#400 value1=32'd502;value2=32'd523;
#400 value1=32'd70;value2=32'd162;
#400 value1=32'd239;value2=32'd253;
#400 value1=32'd306;value2=32'd319;
#400 value1=32'd419;value2=32'd455;
#400 value1=32'd476;value2=32'd477;
#400 value1=32'd484;value2=32'd487;
#400 value1=32'd488;value2=32'd489;
#400 value1=32'd490;value2=32'd491;
#400 value1=32'd527;value2=32'd529;
#400 value1=32'd161;value2=32'd163;
#400 value1=32'd254;value2=32'd305;
#400 value1=32'd307;value2=32'd320;
#400 value1=32'd420;value2=32'd456;
#400 value1=32'd478;value2=32'd483;
#400 value1=32'd487;value2=32'd488;
#400 value1=32'd494;value2=32'd495;
#400 value1=32'd531;value2=32'd533;
#400 value1=32'd164;value2=32'd255;
#400 value1=32'd308;value2=32'd321;
#400 value1=32'd360;value2=32'd421;
#400 value1=32'd441;value2=32'd457;
#400 value1=32'd476;value2=32'd479;
#400 value1=32'd486;value2=32'd487;
#400 value1=32'd494;value2=32'd498;
#400 value1=32'd534;value2=32'd536;
#400 value1=32'd165;value2=32'd256;
#400 value1=32'd309;value2=32'd322;
#400 value1=32'd405;value2=32'd422;
#400 value1=32'd458;value2=32'd476;
#400 value1=32'd480;value2=32'd485;
#400 value1=32'd488;value2=32'd495;
#400 value1=32'd498;value2=32'd538;
#400 value1=32'd166;value2=32'd257;
#400 value1=32'd310;value2=32'd323;
#400 value1=32'd360;value2=32'd423;
#400 value1=32'd441;value2=32'd459;
#400 value1=32'd481;value2=32'd483;
#400 value1=32'd484;value2=32'd485;
#400 value1=32'd488;value2=32'd496;
#400 value1=32'd499;value2=32'd501;
#400 value1=32'd537;value2=32'd539;
#400 value1=32'd167;value2=32'd258;
#400 value1=32'd311;value2=32'd324;
#400 value1=32'd405;value2=32'd424;
#400 value1=32'd460;value2=32'd482;
#400 value1=32'd483;value2=32'd484;
#400 value1=32'd486;value2=32'd487;
#400 value1=32'd497;value2=32'd500;
#400 value1=32'd502;value2=32'd538;
#400 value1=32'd72;value2=32'd162;
#400 value1=32'd241;value2=32'd259;
#400 value1=32'd306;value2=32'd325;
#400 value1=32'd425;value2=32'd461;
#400 value1=32'd478;value2=32'd483;
#400 value1=32'd492;value2=32'd493;
#400 value1=32'd496;value2=32'd497;
#400 value1=32'd541;value2=32'd543;
#400 value1=32'd73;value2=32'd242;
#400 value1=32'd260;value2=32'd326;
#400 value1=32'd361;value2=32'd426;
#400 value1=32'd442;value2=32'd462;
#400 value1=32'd477;value2=32'd479;
#400 value1=32'd483;value2=32'd491;
#400 value1=32'd492;value2=32'd494;
#400 value1=32'd499;value2=32'd500;
#400 value1=32'd544;value2=32'd546;
#400 value1=32'd74;value2=32'd243;
#400 value1=32'd261;value2=32'd327;
#400 value1=32'd406;value2=32'd427;
#400 value1=32'd463;value2=32'd477;
#400 value1=32'd480;value2=32'd483;
#400 value1=32'd490;value2=32'd493;
#400 value1=32'd495;value2=32'd501;
#400 value1=32'd502;value2=32'd548;
#400 value1=32'd75;value2=32'd244;
#400 value1=32'd262;value2=32'd328;
#400 value1=32'd361;value2=32'd428;
#400 value1=32'd442;value2=32'd464;
#400 value1=32'd481;value2=32'd489;
#400 value1=32'd490;value2=32'd493;
#400 value1=32'd496;value2=32'd503;
#400 value1=32'd547;value2=32'd549;
#400 value1=32'd76;value2=32'd245;
#400 value1=32'd263;value2=32'd329;
#400 value1=32'd406;value2=32'd429;
#400 value1=32'd465;value2=32'd482;
#400 value1=32'd489;value2=32'd491;
#400 value1=32'd492;value2=32'd497;
#400 value1=32'd503;value2=32'd548;
#400 value1=32'd164;value2=32'd264;
#400 value1=32'd308;value2=32'd330;
#400 value1=32'd362;value2=32'd430;
#400 value1=32'd443;value2=32'd466;
#400 value1=32'd478;value2=32'd484;
#400 value1=32'd485;value2=32'd490;
#400 value1=32'd495;value2=32'd496;
#400 value1=32'd499;value2=32'd500;
#400 value1=32'd550;value2=32'd552;
#400 value1=32'd165;value2=32'd265;
#400 value1=32'd309;value2=32'd331;
#400 value1=32'd407;value2=32'd431;
#400 value1=32'd467;value2=32'd478;
#400 value1=32'd484;value2=32'd486;
#400 value1=32'd491;value2=32'd494;
#400 value1=32'd497;value2=32'd501;
#400 value1=32'd502;value2=32'd554;
#400 value1=32'd166;value2=32'd266;
#400 value1=32'd310;value2=32'd332;
#400 value1=32'd362;value2=32'd432;
#400 value1=32'd443;value2=32'd468;
#400 value1=32'd487;value2=32'd489;
#400 value1=32'd492;value2=32'd494;
#400 value1=32'd497;value2=32'd503;
#400 value1=32'd553;value2=32'd555;
#400 value1=32'd167;value2=32'd267;
#400 value1=32'd311;value2=32'd333;
#400 value1=32'd407;value2=32'd433;
#400 value1=32'd469;value2=32'd488;
#400 value1=32'd489;value2=32'd493;
#400 value1=32'd495;value2=32'd496;
#400 value1=32'd503;value2=32'd554;
#400 value1=32'd268;value2=32'd334;
#400 value1=32'd364;value2=32'd408;
#400 value1=32'd434;value2=32'd445;
#400 value1=32'd470;value2=32'd479;
#400 value1=32'd480;value2=32'd485;
#400 value1=32'd486;value2=32'd500;
#400 value1=32'd501;value2=32'd557;
#400 value1=32'd269;value2=32'd335;
#400 value1=32'd363;value2=32'd365;
#400 value1=32'd435;value2=32'd444;
#400 value1=32'd446;value2=32'd471;
#400 value1=32'd481;value2=32'd487;
#400 value1=32'd490;value2=32'd494;
#400 value1=32'd500;value2=32'd501;
#400 value1=32'd556;value2=32'd558;
#400 value1=32'd270;value2=32'd336;
#400 value1=32'd366;value2=32'd408;
#400 value1=32'd436;value2=32'd447;
#400 value1=32'd472;value2=32'd482;
#400 value1=32'd488;value2=32'd490;
#400 value1=32'd494;value2=32'd498;
#400 value1=32'd499;value2=32'd502;
#400 value1=32'd503;value2=32'd557;
#400 value1=32'd271;value2=32'd337;
#400 value1=32'd364;value2=32'd410;
#400 value1=32'd437;value2=32'd445;
#400 value1=32'd473;value2=32'd481;
#400 value1=32'd487;value2=32'd491;
#400 value1=32'd495;value2=32'd498;
#400 value1=32'd499;value2=32'd502;
#400 value1=32'd503;value2=32'd559;
#400 value1=32'd272;value2=32'd338;
#400 value1=32'd409;value2=32'd411;
#400 value1=32'd438;value2=32'd474;
#400 value1=32'd482;value2=32'd488;
#400 value1=32'd491;value2=32'd495;
#400 value1=32'd500;value2=32'd501;
#400 value1=32'd273;value2=32'd339;
#400 value1=32'd366;value2=32'd410;
#400 value1=32'd439;value2=32'd447;
#400 value1=32'd475;value2=32'd492;
#400 value1=32'd493;value2=32'd496;
#400 value1=32'd497;value2=32'd500;
#400 value1=32'd501;value2=32'd559;
#400 value1=32'd77;value2=32'd84;
#400 value1=32'd169;value2=32'd246;
#400 value1=32'd253;value2=32'd313;
#400 value1=32'd505;value2=32'd508;
#400 value1=32'd509;value2=32'd510;
#400 value1=32'd511;value2=32'd512;
#400 value1=32'd526;value2=32'd527;
#400 value1=32'd85;value2=32'd168;
#400 value1=32'd170;value2=32'd254;
#400 value1=32'd312;value2=32'd314;
#400 value1=32'd504;value2=32'd508;
#400 value1=32'd509;value2=32'd515;
#400 value1=32'd516;value2=32'd525;
#400 value1=32'd530;value2=32'd531;
#400 value1=32'd86;value2=32'd171;
#400 value1=32'd255;value2=32'd315;
#400 value1=32'd367;value2=32'd448;
#400 value1=32'd507;value2=32'd508;
#400 value1=32'd515;value2=32'd519;
#400 value1=32'd526;value2=32'd534;
#400 value1=32'd87;value2=32'd172;
#400 value1=32'd256;value2=32'd316;
#400 value1=32'd412;value2=32'd476;
#400 value1=32'd506;value2=32'd509;
#400 value1=32'd516;value2=32'd519;
#400 value1=32'd527;value2=32'd534;
#400 value1=32'd88;value2=32'd173;
#400 value1=32'd257;value2=32'd317;
#400 value1=32'd367;value2=32'd448;
#400 value1=32'd504;value2=32'd505;
#400 value1=32'd506;value2=32'd509;
#400 value1=32'd517;value2=32'd520;
#400 value1=32'd522;value2=32'd528;
#400 value1=32'd535;value2=32'd537;
#400 value1=32'd89;value2=32'd174;
#400 value1=32'd258;value2=32'd318;
#400 value1=32'd412;value2=32'd476;
#400 value1=32'd504;value2=32'd505;
#400 value1=32'd507;value2=32'd508;
#400 value1=32'd518;value2=32'd521;
#400 value1=32'd523;value2=32'd529;
#400 value1=32'd536;value2=32'd538;
#400 value1=32'd79;value2=32'd90;
#400 value1=32'd169;value2=32'd248;
#400 value1=32'd259;value2=32'd313;
#400 value1=32'd504;value2=32'd513;
#400 value1=32'd514;value2=32'd517;
#400 value1=32'd518;value2=32'd525;
#400 value1=32'd540;value2=32'd541;
#400 value1=32'd80;value2=32'd91;
#400 value1=32'd249;value2=32'd260;
#400 value1=32'd368;value2=32'd449;
#400 value1=32'd504;value2=32'd512;
#400 value1=32'd513;value2=32'd515;
#400 value1=32'd520;value2=32'd521;
#400 value1=32'd526;value2=32'd544;
#400 value1=32'd81;value2=32'd92;
#400 value1=32'd250;value2=32'd261;
#400 value1=32'd413;value2=32'd477;
#400 value1=32'd504;value2=32'd511;
#400 value1=32'd514;value2=32'd516;
#400 value1=32'd522;value2=32'd523;
#400 value1=32'd527;value2=32'd544;
#400 value1=32'd82;value2=32'd93;
#400 value1=32'd251;value2=32'd262;
#400 value1=32'd368;value2=32'd449;
#400 value1=32'd510;value2=32'd511;
#400 value1=32'd514;value2=32'd517;
#400 value1=32'd524;value2=32'd528;
#400 value1=32'd545;value2=32'd547;
#400 value1=32'd83;value2=32'd94;
#400 value1=32'd252;value2=32'd263;
#400 value1=32'd413;value2=32'd477;
#400 value1=32'd510;value2=32'd512;
#400 value1=32'd513;value2=32'd518;
#400 value1=32'd524;value2=32'd529;
#400 value1=32'd546;value2=32'd548;
#400 value1=32'd95;value2=32'd171;
#400 value1=32'd264;value2=32'd315;
#400 value1=32'd369;value2=32'd450;
#400 value1=32'd505;value2=32'd506;
#400 value1=32'd511;value2=32'd516;
#400 value1=32'd517;value2=32'd520;
#400 value1=32'd521;value2=32'd530;
#400 value1=32'd540;value2=32'd550;
#400 value1=32'd96;value2=32'd172;
#400 value1=32'd265;value2=32'd316;
#400 value1=32'd414;value2=32'd478;
#400 value1=32'd505;value2=32'd507;
#400 value1=32'd512;value2=32'd515;
#400 value1=32'd518;value2=32'd522;
#400 value1=32'd523;value2=32'd531;
#400 value1=32'd541;value2=32'd550;
#400 value1=32'd97;value2=32'd173;
#400 value1=32'd266;value2=32'd317;
#400 value1=32'd369;value2=32'd450;
#400 value1=32'd508;value2=32'd510;
#400 value1=32'd513;value2=32'd515;
#400 value1=32'd518;value2=32'd524;
#400 value1=32'd532;value2=32'd542;
#400 value1=32'd551;value2=32'd553;
#400 value1=32'd98;value2=32'd174;
#400 value1=32'd267;value2=32'd318;
#400 value1=32'd414;value2=32'd478;
#400 value1=32'd509;value2=32'd510;
#400 value1=32'd514;value2=32'd516;
#400 value1=32'd517;value2=32'd524;
#400 value1=32'd533;value2=32'd543;
#400 value1=32'd552;value2=32'd554;
#400 value1=32'd99;value2=32'd268;
#400 value1=32'd371;value2=32'd415;
#400 value1=32'd452;value2=32'd479;
#400 value1=32'd506;value2=32'd507;
#400 value1=32'd521;value2=32'd522;
#400 value1=32'd534;value2=32'd544;
#400 value1=32'd100;value2=32'd269;
#400 value1=32'd370;value2=32'd372;
#400 value1=32'd451;value2=32'd453;
#400 value1=32'd508;value2=32'd511;
#400 value1=32'd515;value2=32'd521;
#400 value1=32'd522;value2=32'd535;
#400 value1=32'd545;value2=32'd556;
#400 value1=32'd101;value2=32'd270;
#400 value1=32'd373;value2=32'd415;
#400 value1=32'd454;value2=32'd479;
#400 value1=32'd509;value2=32'd511;
#400 value1=32'd515;value2=32'd519;
#400 value1=32'd520;value2=32'd523;
#400 value1=32'd524;value2=32'd536;
#400 value1=32'd546;value2=32'd557;
#400 value1=32'd102;value2=32'd271;
#400 value1=32'd371;value2=32'd417;
#400 value1=32'd452;value2=32'd481;
#400 value1=32'd508;value2=32'd512;
#400 value1=32'd516;value2=32'd519;
#400 value1=32'd520;value2=32'd523;
#400 value1=32'd524;value2=32'd537;
#400 value1=32'd547;value2=32'd556;
#400 value1=32'd103;value2=32'd272;
#400 value1=32'd416;value2=32'd418;
#400 value1=32'd480;value2=32'd482;
#400 value1=32'd509;value2=32'd512;
#400 value1=32'd516;value2=32'd521;
#400 value1=32'd522;value2=32'd538;
#400 value1=32'd548;value2=32'd557;
#400 value1=32'd104;value2=32'd273;
#400 value1=32'd373;value2=32'd417;
#400 value1=32'd454;value2=32'd481;
#400 value1=32'd513;value2=32'd514;
#400 value1=32'd517;value2=32'd518;
#400 value1=32'd521;value2=32'd522;
#400 value1=32'd539;value2=32'd549;
#400 value1=32'd558;value2=32'd559;
#400 value1=32'd85;value2=32'd175;
#400 value1=32'd181;value2=32'd254;
#400 value1=32'd319;value2=32'd325;
#400 value1=32'd505;value2=32'd510;
#400 value1=32'd528;value2=32'd529;
#400 value1=32'd532;value2=32'd533;
#400 value1=32'd540;value2=32'd541;
#400 value1=32'd86;value2=32'd182;
#400 value1=32'd255;value2=32'd326;
#400 value1=32'd374;value2=32'd455;
#400 value1=32'd504;value2=32'd506;
#400 value1=32'd511;value2=32'd527;
#400 value1=32'd528;value2=32'd530;
#400 value1=32'd535;value2=32'd536;
#400 value1=32'd540;value2=32'd544;
#400 value1=32'd87;value2=32'd183;
#400 value1=32'd256;value2=32'd327;
#400 value1=32'd419;value2=32'd483;
#400 value1=32'd504;value2=32'd507;
#400 value1=32'd512;value2=32'd526;
#400 value1=32'd529;value2=32'd531;
#400 value1=32'd537;value2=32'd538;
#400 value1=32'd541;value2=32'd544;
#400 value1=32'd88;value2=32'd184;
#400 value1=32'd257;value2=32'd328;
#400 value1=32'd374;value2=32'd455;
#400 value1=32'd508;value2=32'd513;
#400 value1=32'd525;value2=32'd526;
#400 value1=32'd529;value2=32'd532;
#400 value1=32'd539;value2=32'd542;
#400 value1=32'd545;value2=32'd547;
#400 value1=32'd89;value2=32'd185;
#400 value1=32'd258;value2=32'd329;
#400 value1=32'd419;value2=32'd483;
#400 value1=32'd509;value2=32'd514;
#400 value1=32'd525;value2=32'd527;
#400 value1=32'd528;value2=32'd533;
#400 value1=32'd539;value2=32'd543;
#400 value1=32'd546;value2=32'd548;
#400 value1=32'd177;value2=32'd186;
#400 value1=32'd321;value2=32'd330;
#400 value1=32'd375;value2=32'd456;
#400 value1=32'd505;value2=32'd515;
#400 value1=32'd526;value2=32'd531;
#400 value1=32'd532;value2=32'd535;
#400 value1=32'd536;value2=32'd550;
#400 value1=32'd178;value2=32'd187;
#400 value1=32'd322;value2=32'd331;
#400 value1=32'd420;value2=32'd484;
#400 value1=32'd505;value2=32'd516;
#400 value1=32'd527;value2=32'd530;
#400 value1=32'd533;value2=32'd537;
#400 value1=32'd538;value2=32'd550;
#400 value1=32'd179;value2=32'd188;
#400 value1=32'd323;value2=32'd332;
#400 value1=32'd375;value2=32'd456;
#400 value1=32'd517;value2=32'd525;
#400 value1=32'd528;value2=32'd530;
#400 value1=32'd533;value2=32'd539;
#400 value1=32'd551;value2=32'd553;
#400 value1=32'd180;value2=32'd189;
#400 value1=32'd324;value2=32'd333;
#400 value1=32'd420;value2=32'd484;
#400 value1=32'd518;value2=32'd525;
#400 value1=32'd529;value2=32'd531;
#400 value1=32'd532;value2=32'd539;
#400 value1=32'd552;value2=32'd554;
#400 value1=32'd190;value2=32'd334;
#400 value1=32'd377;value2=32'd421;
#400 value1=32'd458;value2=32'd485;
#400 value1=32'd506;value2=32'd507;
#400 value1=32'd519;value2=32'd536;
#400 value1=32'd537;value2=32'd550;
#400 value1=32'd191;value2=32'd335;
#400 value1=32'd376;value2=32'd378;
#400 value1=32'd457;value2=32'd459;
#400 value1=32'd508;value2=32'd520;
#400 value1=32'd526;value2=32'd530;
#400 value1=32'd536;value2=32'd537;
#400 value1=32'd551;value2=32'd556;
#400 value1=32'd192;value2=32'd336;
#400 value1=32'd379;value2=32'd421;
#400 value1=32'd460;value2=32'd485;
#400 value1=32'd509;value2=32'd521;
#400 value1=32'd526;value2=32'd530;
#400 value1=32'd534;value2=32'd535;
#400 value1=32'd538;value2=32'd539;
#400 value1=32'd552;value2=32'd557;
#400 value1=32'd193;value2=32'd337;
#400 value1=32'd377;value2=32'd423;
#400 value1=32'd458;value2=32'd487;
#400 value1=32'd508;value2=32'd522;
#400 value1=32'd527;value2=32'd531;
#400 value1=32'd534;value2=32'd535;
#400 value1=32'd538;value2=32'd539;
#400 value1=32'd553;value2=32'd556;
#400 value1=32'd194;value2=32'd338;
#400 value1=32'd422;value2=32'd424;
#400 value1=32'd486;value2=32'd488;
#400 value1=32'd509;value2=32'd523;
#400 value1=32'd527;value2=32'd531;
#400 value1=32'd536;value2=32'd537;
#400 value1=32'd554;value2=32'd557;
#400 value1=32'd195;value2=32'd339;
#400 value1=32'd379;value2=32'd423;
#400 value1=32'd460;value2=32'd487;
#400 value1=32'd524;value2=32'd528;
#400 value1=32'd529;value2=32'd532;
#400 value1=32'd533;value2=32'd536;
#400 value1=32'd537;value2=32'd555;
#400 value1=32'd558;value2=32'd559;
#400 value1=32'd95;value2=32'd182;
#400 value1=32'd264;value2=32'd326;
#400 value1=32'd380;value2=32'd461;
#400 value1=32'd510;value2=32'd515;
#400 value1=32'd525;value2=32'd526;
#400 value1=32'd541;value2=32'd542;
#400 value1=32'd545;value2=32'd546;
#400 value1=32'd551;value2=32'd552;
#400 value1=32'd96;value2=32'd183;
#400 value1=32'd265;value2=32'd327;
#400 value1=32'd425;value2=32'd489;
#400 value1=32'd510;value2=32'd516;
#400 value1=32'd525;value2=32'd527;
#400 value1=32'd540;value2=32'd543;
#400 value1=32'd547;value2=32'd548;
#400 value1=32'd553;value2=32'd554;
#400 value1=32'd97;value2=32'd184;
#400 value1=32'd266;value2=32'd328;
#400 value1=32'd380;value2=32'd461;
#400 value1=32'd517;value2=32'd528;
#400 value1=32'd540;value2=32'd543;
#400 value1=32'd549;value2=32'd555;
#400 value1=32'd98;value2=32'd185;
#400 value1=32'd267;value2=32'd329;
#400 value1=32'd425;value2=32'd489;
#400 value1=32'd518;value2=32'd529;
#400 value1=32'd541;value2=32'd542;
#400 value1=32'd549;value2=32'd555;
#400 value1=32'd99;value2=32'd268;
#400 value1=32'd382;value2=32'd426;
#400 value1=32'd463;value2=32'd490;
#400 value1=32'd511;value2=32'd512;
#400 value1=32'd519;value2=32'd526;
#400 value1=32'd527;value2=32'd546;
#400 value1=32'd547;value2=32'd550;
#400 value1=32'd556;value2=32'd557;
#400 value1=32'd100;value2=32'd269;
#400 value1=32'd381;value2=32'd383;
#400 value1=32'd462;value2=32'd464;
#400 value1=32'd513;value2=32'd520;
#400 value1=32'd528;value2=32'd540;
#400 value1=32'd546;value2=32'd547;
#400 value1=32'd551;value2=32'd558;
#400 value1=32'd101;value2=32'd270;
#400 value1=32'd384;value2=32'd426;
#400 value1=32'd465;value2=32'd490;
#400 value1=32'd514;value2=32'd521;
#400 value1=32'd529;value2=32'd540;
#400 value1=32'd544;value2=32'd545;
#400 value1=32'd548;value2=32'd549;
#400 value1=32'd552;value2=32'd558;
#400 value1=32'd102;value2=32'd271;
#400 value1=32'd382;value2=32'd428;
#400 value1=32'd463;value2=32'd492;
#400 value1=32'd513;value2=32'd522;
#400 value1=32'd528;value2=32'd541;
#400 value1=32'd544;value2=32'd545;
#400 value1=32'd548;value2=32'd549;
#400 value1=32'd553;value2=32'd559;
#400 value1=32'd103;value2=32'd272;
#400 value1=32'd427;value2=32'd429;
#400 value1=32'd491;value2=32'd493;
#400 value1=32'd514;value2=32'd523;
#400 value1=32'd529;value2=32'd541;
#400 value1=32'd546;value2=32'd547;
#400 value1=32'd554;value2=32'd559;
#400 value1=32'd104;value2=32'd273;
#400 value1=32'd384;value2=32'd428;
#400 value1=32'd465;value2=32'd492;
#400 value1=32'd524;value2=32'd542;
#400 value1=32'd543;value2=32'd546;
#400 value1=32'd547;value2=32'd555;
#400 value1=32'd190;value2=32'd334;
#400 value1=32'd386;value2=32'd430;
#400 value1=32'd467;value2=32'd494;
#400 value1=32'd515;value2=32'd516;
#400 value1=32'd530;value2=32'd531;
#400 value1=32'd534;value2=32'd544;
#400 value1=32'd552;value2=32'd553;
#400 value1=32'd556;value2=32'd557;
#400 value1=32'd191;value2=32'd335;
#400 value1=32'd385;value2=32'd387;
#400 value1=32'd466;value2=32'd468;
#400 value1=32'd517;value2=32'd532;
#400 value1=32'd535;value2=32'd540;
#400 value1=32'd545;value2=32'd552;
#400 value1=32'd553;value2=32'd558;
#400 value1=32'd192;value2=32'd336;
#400 value1=32'd388;value2=32'd430;
#400 value1=32'd469;value2=32'd494;
#400 value1=32'd518;value2=32'd533;
#400 value1=32'd536;value2=32'd540;
#400 value1=32'd546;value2=32'd550;
#400 value1=32'd551;value2=32'd554;
#400 value1=32'd555;value2=32'd558;
#400 value1=32'd193;value2=32'd337;
#400 value1=32'd386;value2=32'd432;
#400 value1=32'd467;value2=32'd496;
#400 value1=32'd517;value2=32'd532;
#400 value1=32'd537;value2=32'd541;
#400 value1=32'd547;value2=32'd550;
#400 value1=32'd551;value2=32'd554;
#400 value1=32'd555;value2=32'd559;
#400 value1=32'd194;value2=32'd338;
#400 value1=32'd431;value2=32'd433;
#400 value1=32'd495;value2=32'd497;
#400 value1=32'd518;value2=32'd533;
#400 value1=32'd538;value2=32'd541;
#400 value1=32'd548;value2=32'd552;
#400 value1=32'd553;value2=32'd559;
#400 value1=32'd195;value2=32'd339;
#400 value1=32'd388;value2=32'd432;
#400 value1=32'd469;value2=32'd496;
#400 value1=32'd539;value2=32'd542;
#400 value1=32'd543;value2=32'd549;
#400 value1=32'd552;value2=32'd553;
#400 value1=32'd389;value2=32'd392;
#400 value1=32'd435;value2=32'd470;
#400 value1=32'd473;value2=32'd499;
#400 value1=32'd520;value2=32'd522;
#400 value1=32'd535;value2=32'd537;
#400 value1=32'd544;value2=32'd550;
#400 value1=32'd557;value2=32'd558;
#400 value1=32'd393;value2=32'd434;
#400 value1=32'd436;value2=32'd474;
#400 value1=32'd498;value2=32'd500;
#400 value1=32'd521;value2=32'd523;
#400 value1=32'd536;value2=32'd538;
#400 value1=32'd544;value2=32'd550;
#400 value1=32'd556;value2=32'd559;
#400 value1=32'd391;value2=32'd394;
#400 value1=32'd435;value2=32'd472;
#400 value1=32'd475;value2=32'd499;
#400 value1=32'd524;value2=32'd539;
#400 value1=32'd545;value2=32'd546;
#400 value1=32'd551;value2=32'd552;
#400 value1=32'd556;value2=32'd559;
#400 value1=32'd393;value2=32'd437;
#400 value1=32'd439;value2=32'd474;
#400 value1=32'd501;value2=32'd503;
#400 value1=32'd524;value2=32'd539;
#400 value1=32'd547;value2=32'd548;
#400 value1=32'd553;value2=32'd554;
#400 value1=32'd557;value2=32'd558;
//rowpointer
#400 value1=8736+1;   value2=8736+14;
#400 value1=8736+28;  value2=8736+40;
#400 value1=8736+52;  value2=8736+68;
#400 value1=8736+84;  value2=8736+98;
#400 value1=8736+112; value2=8736+126;
#400 value1=8736+140; value2=8736+156;
#400 value1=8736+172; value2=8736+188;
#400 value1=8736+204; value2=8736+218;
#400 value1=8736+232; value2=8736+246;
#400 value1=8736+260; value2=8736+274;
#400 value1=8736+286; value2=8736+302;
#400 value1=8736+314; value2=8736+330;
#400 value1=8736+346; value2=8736+362;
#400 value1=8736+378; value2=8736+394;
#400 value1=8736+410; value2=8736+426;
#400 value1=8736+442; value2=8736+458;
#400 value1=8736+474; value2=8736+490;
#400 value1=8736+506; value2=8736+522;
#400 value1=8736+540; value2=8736+558;
#400 value1=8736+576; value2=8736+594;
#400 value1=8736+606; value2=8736+620;
#400 value1=8736+636; value2=8736+650;
#400 value1=8736+666; value2=8736+680;
#400 value1=8736+696; value2=8736+710;
#400 value1=8736+726; value2=8736+740;
#400 value1=8736+756; value2=8736+772;
#400 value1=8736+786; value2=8736+800;
#400 value1=8736+816; value2=8736+830;
#400 value1=8736+846; value2=8736+862;
#400 value1=8736+876; value2=8736+892;
#400 value1=8736+906; value2=8736+922;
#400 value1=8736+938; value2=8736+956;
#400 value1=8736+972; value2=8736+990;
#400 value1=8736+1006;value2=8736+1024;
#400 value1=8736+1040;value2=8736+1058;
#400 value1=8736+1074;value2=8736+1092;
#400 value1=8736+1108;value2=8736+1126;
#400 value1=8736+1144;value2=8736+1160;
#400 value1=8736+1178;value2=8736+1194;
#400 value1=8736+1208;value2=8736+1220;
#400 value1=8736+1236;value2=8736+1250;
#400 value1=8736+1264;value2=8736+1280;
#400 value1=8736+1296;value2=8736+1312;
#400 value1=8736+1328;value2=8736+1344;
#400 value1=8736+1360;value2=8736+1378;
#400 value1=8736+1396;value2=8736+1410;
#400 value1=8736+1426;value2=8736+1442;
#400 value1=8736+1456;value2=8736+1470;
#400 value1=8736+1488;value2=8736+1506;
#400 value1=8736+1522;value2=8736+1538;
#400 value1=8736+1554;value2=8736+1570;
#400 value1=8736+1588;value2=8736+1606;
#400 value1=8736+1622;value2=8736+1638;
#400 value1=8736+1652;value2=8736+1668;
#400 value1=8736+1684;value2=8736+1700;
#400 value1=8736+1716;value2=8736+1732;
#400 value1=8736+1748;value2=8736+1764;
#400 value1=8736+1780;value2=8736+1798;
#400 value1=8736+1816;value2=8736+1834;
#400 value1=8736+1852;value2=8736+1866;
#400 value1=8736+1880;value2=8736+1894;
#400 value1=8736+1908;value2=8736+1924;
#400 value1=8736+1936;value2=8736+1952;
#400 value1=8736+1964;value2=8736+1980;
#400 value1=8736+1996;value2=8736+2012;
#400 value1=8736+2028;value2=8736+2040;
#400 value1=8736+2054;value2=8736+2070;
#400 value1=8736+2086;value2=8736+2100;
#400 value1=8736+2116;value2=8736+2130;
#400 value1=8736+2144;value2=8736+2160;
#400 value1=8736+2174;value2=8736+2190;
#400 value1=8736+2206;value2=8736+2220;
#400 value1=8736+2236;value2=8736+2250;
#400 value1=8736+2266;value2=8736+2280;
#400 value1=8736+2296;value2=8736+2310;
#400 value1=8736+2326;value2=8736+2340;
#400 value1=8736+2356;value2=8736+2374;
#400 value1=8736+2390;value2=8736+2408;
#400 value1=8736+2424;value2=8736+2440;
#400 value1=8736+2458;value2=8736+2474;
#400 value1=8736+2492;value2=8736+2510;
#400 value1=8736+2526;value2=8736+2544;
#400 value1=8736+2560;value2=8736+2578;
#400 value1=8736+2594;value2=8736+2612;
#400 value1=8736+2628;value2=8736+2642;
#400 value1=8736+2658;value2=8736+2674;
#400 value1=8736+2690;value2=8736+2706;
#400 value1=8736+2724;value2=8736+2742;
#400 value1=8736+2758;value2=8736+2770;
#400 value1=8736+2784;value2=8736+2798;
#400 value1=8736+2814;value2=8736+2830;
#400 value1=8736+2844;value2=8736+2862;
#400 value1=8736+2880;value2=8736+2896;
#400 value1=8736+2912;value2=8736+2928;
#400 value1=8736+2944;value2=8736+2958;
#400 value1=8736+2972;value2=8736+2988;
#400 value1=8736+3004;value2=8736+3022;
#400 value1=8736+3040;value2=8736+3056;
#400 value1=8736+3072;value2=8736+3088;
#400 value1=8736+3104;value2=8736+3116;
#400 value1=8736+3128;value2=8736+3142;
#400 value1=8736+3156;value2=8736+3170;
#400 value1=8736+3184;value2=8736+3200;
#400 value1=8736+3216;value2=8736+3232;
#400 value1=8736+3248;value2=8736+3264;
#400 value1=8736+3278;value2=8736+3294;
#400 value1=8736+3310;value2=8736+3328;
#400 value1=8736+3344;value2=8736+3362;
#400 value1=8736+3378;value2=8736+3396;
#400 value1=8736+3412;value2=8736+3430;
#400 value1=8736+3446;value2=8736+3460;
#400 value1=8736+3476;value2=8736+3494;
#400 value1=8736+3510;value2=8736+3528;
#400 value1=8736+3546;value2=8736+3562;
#400 value1=8736+3580;value2=8736+3596;
#400 value1=8736+3608;value2=8736+3622;
#400 value1=8736+3638;value2=8736+3652;
#400 value1=8736+3668;value2=8736+3682;
#400 value1=8736+3698;value2=8736+3712;
#400 value1=8736+3728;value2=8736+3742;
#400 value1=8736+3758;value2=8736+3772;
#400 value1=8736+3788;value2=8736+3804;
#400 value1=8736+3818;value2=8736+3834;
#400 value1=8736+3848;value2=8736+3862;
#400 value1=8736+3874;value2=8736+3890;
#400 value1=8736+3904;value2=8736+3918;
#400 value1=8736+3934;value2=8736+3950;
#400 value1=8736+3966;value2=8736+3982;
#400 value1=8736+3998;value2=8736+4014;
#400 value1=8736+4032;value2=8736+4050;
#400 value1=8736+4064;value2=8736+4080;
#400 value1=8736+4096;value2=8736+4110;
#400 value1=8736+4124;value2=8736+4142;
#400 value1=8736+4160;value2=8736+4176;
#400 value1=8736+4192;value2=8736+4208;
#400 value1=8736+4224;value2=8736+4242;
#400 value1=8736+4260;value2=8736+4276;
#400 value1=8736+4292;value2=8736+4308;
#400 value1=8736+4322;value2=8736+4338;
#400 value1=8736+4356;value2=8736+4372;
#400 value1=8736+4390;value2=8736+4406;
#400 value1=8736+4422;value2=8736+4440;
#400 value1=8736+4456;value2=8736+4474;
#400 value1=8736+4490;value2=8736+4504;
#400 value1=8736+4522;value2=8736+4538;
#400 value1=8736+4556;value2=8736+4572;
#400 value1=8736+4590;value2=8736+4606;
#400 value1=8736+4624;value2=8736+4640;
#400 value1=8736+4652;value2=8736+4668;
#400 value1=8736+4682;value2=8736+4698;
#400 value1=8736+4712;value2=8736+4726;
#400 value1=8736+4742;value2=8736+4756;
#400 value1=8736+4772;value2=8736+4788;
#400 value1=8736+4802;value2=8736+4818;
#400 value1=8736+4832;value2=8736+4848;
#400 value1=8736+4862;value2=8736+4878;
#400 value1=8736+4892;value2=8736+4906;
#400 value1=8736+4922;value2=8736+4938;
#400 value1=8736+4954;value2=8736+4970;
#400 value1=8736+4988;value2=8736+5006;
#400 value1=8736+5022;value2=8736+5034;
#400 value1=8736+5048;value2=8736+5062;
#400 value1=8736+5078;value2=8736+5094;
#400 value1=8736+5108;value2=8736+5126;
#400 value1=8736+5144;value2=8736+5160;
#400 value1=8736+5176;value2=8736+5192;
#400 value1=8736+5208;value2=8736+5222;
#400 value1=8736+5236;value2=8736+5252;
#400 value1=8736+5268;value2=8736+5286;
#400 value1=8736+5304;value2=8736+5320;
#400 value1=8736+5336;value2=8736+5350;
#400 value1=8736+5364;value2=8736+5380;
#400 value1=8736+5396;value2=8736+5412;
#400 value1=8736+5428;value2=8736+5442;
#400 value1=8736+5456;value2=8736+5470;
#400 value1=8736+5484;value2=8736+5498;
#400 value1=8736+5514;value2=8736+5530;
#400 value1=8736+5546;value2=8736+5562;
#400 value1=8736+5574;value2=8736+5590;
#400 value1=8736+5602;value2=8736+5618;
#400 value1=8736+5636;value2=8736+5654;
#400 value1=8736+5672;value2=8736+5690;
#400 value1=8736+5706;value2=8736+5722;
#400 value1=8736+5738;value2=8736+5754;
#400 value1=8736+5770;value2=8736+5786;
#400 value1=8736+5804;value2=8736+5818;
#400 value1=8736+5834;value2=8736+5850;
#400 value1=8736+5868;value2=8736+5886;
#400 value1=8736+5902;value2=8736+5916;
#400 value1=8736+5932;value2=8736+5948;
#400 value1=8736+5966;value2=8736+5982;
#400 value1=8736+5998;value2=8736+6016;
#400 value1=8736+6030;value2=8736+6046;
#400 value1=8736+6062;value2=8736+6080;
#400 value1=8736+6094;value2=8736+6110;
#400 value1=8736+6124;value2=8736+6136;
#400 value1=8736+6152;value2=8736+6168;
#400 value1=8736+6184;value2=8736+6198;
#400 value1=8736+6212;value2=8736+6230;
#400 value1=8736+6248;value2=8736+6266;
#400 value1=8736+6284;value2=8736+6300;
#400 value1=8736+6316;value2=8736+6332;
#400 value1=8736+6348;value2=8736+6364;
#400 value1=8736+6380;value2=8736+6396;
#400 value1=8736+6412;value2=8736+6428;
#400 value1=8736+6440;value2=8736+6456;
#400 value1=8736+6468;value2=8736+6484;
#400 value1=8736+6500;value2=8736+6518;
#400 value1=8736+6534;value2=8736+6548;
#400 value1=8736+6566;value2=8736+6582;
#400 value1=8736+6600;value2=8736+6616;
#400 value1=8736+6632;value2=8736+6646;
#400 value1=8736+6664;value2=8736+6680;
#400 value1=8736+6696;value2=8736+6714;
#400 value1=8736+6730;value2=8736+6746;
#400 value1=8736+6760;value2=8736+6778;
#400 value1=8736+6794;value2=8736+6810;
#400 value1=8736+6824;value2=8736+6838;
#400 value1=8736+6854;value2=8736+6870;
#400 value1=8736+6886;value2=8736+6898;
#400 value1=8736+6912;value2=8736+6928;
#400 value1=8736+6944;value2=8736+6960;
#400 value1=8736+6976;value2=8736+6990;
#400 value1=8736+7004;value2=8736+7018;
#400 value1=8736+7032;value2=8736+7048;
#400 value1=8736+7064;value2=8736+7082;
#400 value1=8736+7096;value2=8736+7112;
#400 value1=8736+7128;value2=8736+7146;
#400 value1=8736+7164;value2=8736+7180;
#400 value1=8736+7194;value2=8736+7210;
#400 value1=8736+7226;value2=8736+7244;
#400 value1=8736+7260;value2=8736+7276;
#400 value1=8736+7294;value2=8736+7308;
#400 value1=8736+7324;value2=8736+7340;
#400 value1=8736+7358;value2=8736+7372;
#400 value1=8736+7388;value2=8736+7402;
#400 value1=8736+7414;value2=8736+7430;
#400 value1=8736+7446;value2=8736+7462;
#400 value1=8736+7476;value2=8736+7492;
#400 value1=8736+7508;value2=8736+7526;
#400 value1=8736+7542;value2=8736+7556;
#400 value1=8736+7574;value2=8736+7590;
#400 value1=8736+7608;value2=8736+7624;
#400 value1=8736+7640;value2=8736+7654;
#400 value1=8736+7672;value2=8736+7688;
#400 value1=8736+7704;value2=8736+7722;
#400 value1=8736+7738;value2=8736+7754;
#400 value1=8736+7768;value2=8736+7786;
#400 value1=8736+7802;value2=8736+7818;
#400 value1=8736+7832;value2=8736+7846;
#400 value1=8736+7862;value2=8736+7878;
#400 value1=8736+7894;value2=8736+7906;
#400 value1=8736+7920;value2=8736+7934;
#400 value1=8736+7948;value2=8736+7960;
#400 value1=8736+7972;value2=8736+7988;
#400 value1=8736+8004;value2=8736+8018;
#400 value1=8736+8032;value2=8736+8046;
#400 value1=8736+8060;value2=8736+8074;
#400 value1=8736+8090;value2=8736+8106;
#400 value1=8736+8122;value2=8736+8138;
#400 value1=8736+8150;value2=8736+8164;
#400 value1=8736+8180;value2=8736+8196;
#400 value1=8736+8210;value2=8736+8226;
#400 value1=8736+8240;value2=8736+8256;
#400 value1=8736+8272;value2=8736+8288;
#400 value1=8736+8304;value2=8736+8318;
#400 value1=8736+8332;value2=8736+8346;
#400 value1=8736+8360;value2=8736+8372;
#400 value1=8736+8386;value2=8736+8402;
#400 value1=8736+8418;value2=8736+8432;
#400 value1=8736+8448;value2=8736+8464;
#400 value1=8736+8480;value2=8736+8492;
#400 value1=8736+8504;value2=8736+8520;
#400 value1=8736+8534;value2=8736+8550;
#400 value1=8736+8566;value2=8736+8580;
#400 value1=8736+8592;value2=8736+8608;
#400 value1=8736+8622;value2=8736+8638;
#400 value1=8736+8654;value2=8736+8668;
#400 value1=8736+8680;value2=8736+8694;
#400 value1=8736+8708;value2=8736+8722;
#400 value1=8736+8736;value2=0;
//end


//initial begin
#700 value1=0;value2=1;
#400 value1=2;value2=3;
#400 value1=4;value2=5;
#400 value1=6;value2=7;
#400 value1=8;value2=9;
#400 value1=10;value2=11;
#400 value1=12;value2=13;
#400 value1=14;value2=15;
#400 value1=16;value2=17;
#400 value1=18;value2=19;
#400 value1=20;value2=21;
#400 value1=22;value2=23;
#400 value1=24;value2=25;
#400 value1=26;value2=27;
#400 value1=28;value2=29;
#400 value1=30;value2=31;
#400 value1=32;value2=33;
#400 value1=34;value2=35;
#400 value1=36;value2=37;
#400 value1=38;value2=39;
#400 value1=40;value2=41;
#400 value1=42;value2=43;
#400 value1=44;value2=45;
#400 value1=46;value2=47;
#400 value1=48;value2=49;
#400 value1=50;value2=51;
#400 value1=52;value2=53;
#400 value1=54;value2=55;
#400 value1=56;value2=57;
#400 value1=58;value2=59;
#400 value1=60;value2=61;
#400 value1=62;value2=63;
#400 value1=64;value2=65;
#400 value1=66;value2=67;
#400 value1=68;value2=69;
#400 value1=70;value2=71;
#400 value1=72;value2=73;
#400 value1=74;value2=75;
#400 value1=76;value2=77;
#400 value1=78;value2=79;
#400 value1=80;value2=81;
#400 value1=82;value2=83;
#400 value1=84;value2=85;
#400 value1=86;value2=87;
#400 value1=88;value2=89;
#400 value1=90;value2=91;
#400 value1=92;value2=93;
#400 value1=94;value2=95;
#400 value1=96;value2=97;
#400 value1=98;value2=99;
#400 value1=100;value2=101;
#400 value1=102;value2=103;
#400 value1=104;value2=105;
#400 value1=106;value2=107;
#400 value1=108;value2=109;
#400 value1=110;value2=111;
#400 value1=112;value2=113;
#400 value1=114;value2=115;
#400 value1=116;value2=117;
#400 value1=118;value2=119;
#400 value1=120;value2=121;
#400 value1=122;value2=123;
#400 value1=124;value2=125;
#400 value1=126;value2=127;
#400 value1=128;value2=129;
#400 value1=130;value2=131;
#400 value1=132;value2=133;
#400 value1=134;value2=135;
#400 value1=136;value2=137;
#400 value1=138;value2=139;
#400 value1=140;value2=141;
#400 value1=142;value2=143;
#400 value1=144;value2=145;
#400 value1=146;value2=147;
#400 value1=148;value2=149;
#400 value1=150;value2=151;
#400 value1=152;value2=153;
#400 value1=154;value2=155;
#400 value1=156;value2=157;
#400 value1=158;value2=159;
#400 value1=160;value2=161;
#400 value1=162;value2=163;
#400 value1=164;value2=165;
#400 value1=166;value2=167;
#400 value1=168;value2=169;
#400 value1=170;value2=171;
#400 value1=172;value2=173;
#400 value1=174;value2=175;
#400 value1=176;value2=177;
#400 value1=178;value2=179;
#400 value1=180;value2=181;
#400 value1=182;value2=183;
#400 value1=184;value2=185;
#400 value1=186;value2=187;
#400 value1=188;value2=189;
#400 value1=190;value2=191;
#400 value1=192;value2=193;
#400 value1=194;value2=195;
#400 value1=196;value2=197;
#400 value1=198;value2=199;
#400 value1=200;value2=201;
#400 value1=202;value2=203;
#400 value1=204;value2=205;
#400 value1=206;value2=207;
#400 value1=208;value2=209;
#400 value1=210;value2=211;
#400 value1=212;value2=213;
#400 value1=214;value2=215;
#400 value1=216;value2=217;
#400 value1=218;value2=219;
#400 value1=220;value2=221;
#400 value1=222;value2=223;
#400 value1=224;value2=225;
#400 value1=226;value2=227;
#400 value1=228;value2=229;
#400 value1=230;value2=231;
#400 value1=232;value2=233;
#400 value1=234;value2=235;
#400 value1=236;value2=237;
#400 value1=238;value2=239;
#400 value1=240;value2=241;
#400 value1=242;value2=243;
#400 value1=244;value2=245;
#400 value1=246;value2=247;
#400 value1=248;value2=249;
#400 value1=250;value2=251;
#400 value1=252;value2=253;
#400 value1=254;value2=255;
#400 value1=256;value2=257;
#400 value1=258;value2=259;
#400 value1=260;value2=261;
#400 value1=262;value2=263;
#400 value1=264;value2=265;
#400 value1=266;value2=267;
#400 value1=268;value2=269;
#400 value1=270;value2=271;
#400 value1=272;value2=273;
#400 value1=274;value2=275;
#400 value1=276;value2=277;
#400 value1=278;value2=279;
#400 value1=280;value2=281;
#400 value1=282;value2=283;
#400 value1=284;value2=285;
#400 value1=286;value2=287;
#400 value1=288;value2=289;
#400 value1=290;value2=291;
#400 value1=292;value2=293;
#400 value1=294;value2=295;
#400 value1=296;value2=297;
#400 value1=298;value2=299;
#400 value1=300;value2=301;
#400 value1=302;value2=303;
#400 value1=304;value2=305;
#400 value1=306;value2=307;
#400 value1=308;value2=309;
#400 value1=310;value2=311;
#400 value1=312;value2=313;
#400 value1=314;value2=315;
#400 value1=316;value2=317;
#400 value1=318;value2=319;
#400 value1=320;value2=321;
#400 value1=322;value2=323;
#400 value1=324;value2=325;
#400 value1=326;value2=327;
#400 value1=328;value2=329;
#400 value1=330;value2=331;
#400 value1=332;value2=333;
#400 value1=334;value2=335;
#400 value1=336;value2=337;
#400 value1=338;value2=339;
#400 value1=340;value2=341;
#400 value1=342;value2=343;
#400 value1=344;value2=345;
#400 value1=346;value2=347;
#400 value1=348;value2=349;
#400 value1=350;value2=351;
#400 value1=352;value2=353;
#400 value1=354;value2=355;
#400 value1=356;value2=357;
#400 value1=358;value2=359;
#400 value1=360;value2=361;
#400 value1=362;value2=363;
#400 value1=364;value2=365;
#400 value1=366;value2=367;
#400 value1=368;value2=369;
#400 value1=370;value2=371;
#400 value1=372;value2=373;
#400 value1=374;value2=375;
#400 value1=376;value2=377;
#400 value1=378;value2=379;
#400 value1=380;value2=381;
#400 value1=382;value2=383;
#400 value1=384;value2=385;
#400 value1=386;value2=387;
#400 value1=388;value2=389;
#400 value1=390;value2=391;
#400 value1=392;value2=393;
#400 value1=394;value2=395;
#400 value1=396;value2=397;
#400 value1=398;value2=399;
#400 value1=400;value2=401;
#400 value1=402;value2=403;
#400 value1=404;value2=405;
#400 value1=406;value2=407;
#400 value1=408;value2=409;
#400 value1=410;value2=411;
#400 value1=412;value2=413;
#400 value1=414;value2=415;
#400 value1=416;value2=417;
#400 value1=418;value2=419;
#400 value1=420;value2=421;
#400 value1=422;value2=423;
#400 value1=424;value2=425;
#400 value1=426;value2=427;
#400 value1=428;value2=429;
#400 value1=430;value2=431;
#400 value1=432;value2=433;
#400 value1=434;value2=435;
#400 value1=436;value2=437;
#400 value1=438;value2=439;
#400 value1=440;value2=441;
#400 value1=442;value2=443;
#400 value1=444;value2=445;
#400 value1=446;value2=447;
#400 value1=448;value2=449;
#400 value1=450;value2=451;
#400 value1=452;value2=453;
#400 value1=454;value2=455;
#400 value1=456;value2=457;
#400 value1=458;value2=459;
#400 value1=460;value2=461;
#400 value1=462;value2=463;
#400 value1=464;value2=465;
#400 value1=466;value2=467;
#400 value1=468;value2=469;
#400 value1=470;value2=471;
#400 value1=472;value2=473;
#400 value1=474;value2=475;
#400 value1=476;value2=477;
#400 value1=478;value2=479;
#400 value1=480;value2=481;
#400 value1=482;value2=483;
#400 value1=484;value2=485;
#400 value1=486;value2=487;
#400 value1=488;value2=489;
#400 value1=490;value2=491;
#400 value1=492;value2=493;
#400 value1=494;value2=495;
#400 value1=496;value2=497;
#400 value1=498;value2=499;
#400 value1=500;value2=501;
#400 value1=502;value2=503;
#400 value1=504;value2=505;
#400 value1=506;value2=507;
#400 value1=508;value2=509;
#400 value1=510;value2=511;
#400 value1=512;value2=513;
#400 value1=514;value2=515;
#400 value1=516;value2=517;
#400 value1=518;value2=519;
#400 value1=520;value2=521;
#400 value1=522;value2=523;
#400 value1=524;value2=525;
#400 value1=526;value2=527;
#400 value1=528;value2=529;
#400 value1=530;value2=531;
#400 value1=532;value2=533;
#400 value1=534;value2=535;
#400 value1=536;value2=537;
#400 value1=538;value2=539;
#400 value1=540;value2=541;
#400 value1=542;value2=543;
#400 value1=544;value2=545;
#400 value1=546;value2=547;
#400 value1=548;value2=549;
#400 value1=550;value2=551;
#400 value1=552;value2=553;
#400 value1=554;value2=555;
#400 value1=556;value2=557;
#400 value1=558;value2=559;

#34 value1=0;value2=1;
#400 value1=2;value2=3;
#400 value1=4;value2=5;
#400 value1=6;value2=7;
#400 value1=8;value2=9;
#400 value1=10;value2=11;
#400 value1=12;value2=13;
#400 value1=14;value2=15;
#400 value1=16;value2=17;
#400 value1=18;value2=19;
#400 value1=20;value2=21;
#400 value1=22;value2=23;
#400 value1=24;value2=25;
#400 value1=26;value2=27;
#400 value1=28;value2=29;
#400 value1=30;value2=31;
#400 value1=32;value2=33;
#400 value1=34;value2=35;
#400 value1=36;value2=37;
#400 value1=38;value2=39;
#400 value1=40;value2=41;
#400 value1=42;value2=43;
#400 value1=44;value2=45;
#400 value1=46;value2=47;
#400 value1=48;value2=49;
#400 value1=50;value2=51;
#400 value1=52;value2=53;
#400 value1=54;value2=55;
#400 value1=56;value2=57;
#400 value1=58;value2=59;
#400 value1=60;value2=61;
#400 value1=62;value2=63;
#400 value1=64;value2=65;
#400 value1=66;value2=67;
#400 value1=68;value2=69;
#400 value1=70;value2=71;
#400 value1=72;value2=73;
#400 value1=74;value2=75;
#400 value1=76;value2=77;
#400 value1=78;value2=79;
#400 value1=80;value2=81;
#400 value1=82;value2=83;
#400 value1=84;value2=85;
#400 value1=86;value2=87;
#400 value1=88;value2=89;
#400 value1=90;value2=91;
#400 value1=92;value2=93;
#400 value1=94;value2=95;
#400 value1=96;value2=97;
#400 value1=98;value2=99;
#400 value1=100;value2=101;
#400 value1=102;value2=103;
#400 value1=104;value2=105;
#400 value1=106;value2=107;
#400 value1=108;value2=109;
#400 value1=110;value2=111;
#400 value1=112;value2=113;
#400 value1=114;value2=115;
#400 value1=116;value2=117;
#400 value1=118;value2=119;
#400 value1=120;value2=121;
#400 value1=122;value2=123;
#400 value1=124;value2=125;
#400 value1=126;value2=127;
#400 value1=128;value2=129;
#400 value1=130;value2=131;
#400 value1=132;value2=133;
#400 value1=134;value2=135;
#400 value1=136;value2=137;
#400 value1=138;value2=139;
#400 value1=140;value2=141;
#400 value1=142;value2=143;
#400 value1=144;value2=145;
#400 value1=146;value2=147;
#400 value1=148;value2=149;
#400 value1=150;value2=151;
#400 value1=152;value2=153;
#400 value1=154;value2=155;
#400 value1=156;value2=157;
#400 value1=158;value2=159;
#400 value1=160;value2=161;
#400 value1=162;value2=163;
#400 value1=164;value2=165;
#400 value1=166;value2=167;
#400 value1=168;value2=169;
#400 value1=170;value2=171;
#400 value1=172;value2=173;
#400 value1=174;value2=175;
#400 value1=176;value2=177;
#400 value1=178;value2=179;
#400 value1=180;value2=181;
#400 value1=182;value2=183;
#400 value1=184;value2=185;
#400 value1=186;value2=187;
#400 value1=188;value2=189;
#400 value1=190;value2=191;
#400 value1=192;value2=193;
#400 value1=194;value2=195;
#400 value1=196;value2=197;
#400 value1=198;value2=199;
#400 value1=200;value2=201;
#400 value1=202;value2=203;
#400 value1=204;value2=205;
#400 value1=206;value2=207;
#400 value1=208;value2=209;
#400 value1=210;value2=211;
#400 value1=212;value2=213;
#400 value1=214;value2=215;
#400 value1=216;value2=217;
#400 value1=218;value2=219;
#400 value1=220;value2=221;
#400 value1=222;value2=223;
#400 value1=224;value2=225;
#400 value1=226;value2=227;
#400 value1=228;value2=229;
#400 value1=230;value2=231;
#400 value1=232;value2=233;
#400 value1=234;value2=235;
#400 value1=236;value2=237;
#400 value1=238;value2=239;
#400 value1=240;value2=241;
#400 value1=242;value2=243;
#400 value1=244;value2=245;
#400 value1=246;value2=247;
#400 value1=248;value2=249;
#400 value1=250;value2=251;
#400 value1=252;value2=253;
#400 value1=254;value2=255;
#400 value1=256;value2=257;
#400 value1=258;value2=259;
#400 value1=260;value2=261;
#400 value1=262;value2=263;
#400 value1=264;value2=265;
#400 value1=266;value2=267;
#400 value1=268;value2=269;
#400 value1=270;value2=271;
#400 value1=272;value2=273;
#400 value1=274;value2=275;
#400 value1=276;value2=277;
#400 value1=278;value2=279;
#400 value1=280;value2=281;
#400 value1=282;value2=283;
#400 value1=284;value2=285;
#400 value1=286;value2=287;
#400 value1=288;value2=289;
#400 value1=290;value2=291;
#400 value1=292;value2=293;
#400 value1=294;value2=295;
#400 value1=296;value2=297;
#400 value1=298;value2=299;
#400 value1=300;value2=301;
#400 value1=302;value2=303;
#400 value1=304;value2=305;
#400 value1=306;value2=307;
#400 value1=308;value2=309;
#400 value1=310;value2=311;
#400 value1=312;value2=313;
#400 value1=314;value2=315;
#400 value1=316;value2=317;
#400 value1=318;value2=319;
#400 value1=320;value2=321;
#400 value1=322;value2=323;
#400 value1=324;value2=325;
#400 value1=326;value2=327;
#400 value1=328;value2=329;
#400 value1=330;value2=331;
#400 value1=332;value2=333;
#400 value1=334;value2=335;
#400 value1=336;value2=337;
#400 value1=338;value2=339;
#400 value1=340;value2=341;
#400 value1=342;value2=343;
#400 value1=344;value2=345;
#400 value1=346;value2=347;
#400 value1=348;value2=349;
#400 value1=350;value2=351;
#400 value1=352;value2=353;
#400 value1=354;value2=355;
#400 value1=356;value2=357;
#400 value1=358;value2=359;
#400 value1=360;value2=361;
#400 value1=362;value2=363;
#400 value1=364;value2=365;
#400 value1=366;value2=367;
#400 value1=368;value2=369;
#400 value1=370;value2=371;
#400 value1=372;value2=373;
#400 value1=374;value2=375;
#400 value1=376;value2=377;
#400 value1=378;value2=379;
#400 value1=380;value2=381;
#400 value1=382;value2=383;
#400 value1=384;value2=385;
#400 value1=386;value2=387;
#400 value1=388;value2=389;
#400 value1=390;value2=391;
#400 value1=392;value2=393;
#400 value1=394;value2=395;
#400 value1=396;value2=397;
#400 value1=398;value2=399;
#400 value1=400;value2=401;
#400 value1=402;value2=403;
#400 value1=404;value2=405;
#400 value1=406;value2=407;
#400 value1=408;value2=409;
#400 value1=410;value2=411;
#400 value1=412;value2=413;
#400 value1=414;value2=415;
#400 value1=416;value2=417;
#400 value1=418;value2=419;
#400 value1=420;value2=421;
#400 value1=422;value2=423;
#400 value1=424;value2=425;
#400 value1=426;value2=427;
#400 value1=428;value2=429;
#400 value1=430;value2=431;
#400 value1=432;value2=433;
#400 value1=434;value2=435;
#400 value1=436;value2=437;
#400 value1=438;value2=439;
#400 value1=440;value2=441;
#400 value1=442;value2=443;
#400 value1=444;value2=445;
#400 value1=446;value2=447;
#400 value1=448;value2=449;
#400 value1=450;value2=451;
#400 value1=452;value2=453;
#400 value1=454;value2=455;
#400 value1=456;value2=457;
#400 value1=458;value2=459;
#400 value1=460;value2=461;
#400 value1=462;value2=463;
#400 value1=464;value2=465;
#400 value1=466;value2=467;
#400 value1=468;value2=469;
#400 value1=470;value2=471;
#400 value1=472;value2=473;
#400 value1=474;value2=475;
#400 value1=476;value2=477;
#400 value1=478;value2=479;
#400 value1=480;value2=481;
#400 value1=482;value2=483;
#400 value1=484;value2=485;
#400 value1=486;value2=487;
#400 value1=488;value2=489;
#400 value1=490;value2=491;
#400 value1=492;value2=493;
#400 value1=494;value2=495;
#400 value1=496;value2=497;
#400 value1=498;value2=499;
#400 value1=500;value2=501;
#400 value1=502;value2=503;
#400 value1=504;value2=505;
#400 value1=506;value2=507;
#400 value1=508;value2=509;
#400 value1=510;value2=511;
#400 value1=512;value2=513;
#400 value1=514;value2=515;
#400 value1=516;value2=517;
#400 value1=518;value2=519;
#400 value1=520;value2=521;
#400 value1=522;value2=523;
#400 value1=524;value2=525;
#400 value1=526;value2=527;
#400 value1=528;value2=529;
#400 value1=530;value2=531;
#400 value1=532;value2=533;
#400 value1=534;value2=535;
#400 value1=536;value2=537;
#400 value1=538;value2=539;
#400 value1=540;value2=541;
#400 value1=542;value2=543;
#400 value1=544;value2=545;
#400 value1=546;value2=547;
#400 value1=548;value2=549;
#400 value1=550;value2=551;
#400 value1=552;value2=553;
#400 value1=554;value2=555;
#400 value1=556;value2=557;
#400 value1=558;value2=559;
end


endmodule
